module gw_gao(
    \CSI2RAW8_inst/burst_done ,
    \CSI2RAW8_inst/hs_en ,
    \CSI2RAW8_inst/term_en ,
    \CSI2RAW8_inst/lv_8bit ,
    \CSI2RAW8_inst/data[15] ,
    \CSI2RAW8_inst/data[14] ,
    \CSI2RAW8_inst/data[13] ,
    \CSI2RAW8_inst/data[12] ,
    \CSI2RAW8_inst/data[11] ,
    \CSI2RAW8_inst/data[10] ,
    \CSI2RAW8_inst/data[9] ,
    \CSI2RAW8_inst/data[8] ,
    \CSI2RAW8_inst/data[7] ,
    \CSI2RAW8_inst/data[6] ,
    \CSI2RAW8_inst/data[5] ,
    \CSI2RAW8_inst/data[4] ,
    \CSI2RAW8_inst/data[3] ,
    \CSI2RAW8_inst/data[2] ,
    \CSI2RAW8_inst/data[1] ,
    \CSI2RAW8_inst/data[0] ,
    \CSI2RAW8_inst/u_control_capture/cnt[15] ,
    \CSI2RAW8_inst/u_control_capture/cnt[14] ,
    \CSI2RAW8_inst/u_control_capture/cnt[13] ,
    \CSI2RAW8_inst/u_control_capture/cnt[12] ,
    \CSI2RAW8_inst/u_control_capture/cnt[11] ,
    \CSI2RAW8_inst/u_control_capture/cnt[10] ,
    \CSI2RAW8_inst/u_control_capture/cnt[9] ,
    \CSI2RAW8_inst/u_control_capture/cnt[8] ,
    \CSI2RAW8_inst/u_control_capture/cnt[7] ,
    \CSI2RAW8_inst/u_control_capture/cnt[6] ,
    \CSI2RAW8_inst/u_control_capture/cnt[5] ,
    \CSI2RAW8_inst/u_control_capture/cnt[4] ,
    \CSI2RAW8_inst/u_control_capture/cnt[3] ,
    \CSI2RAW8_inst/u_control_capture/cnt[2] ,
    \CSI2RAW8_inst/u_control_capture/cnt[1] ,
    \CSI2RAW8_inst/u_control_capture/cnt[0] ,
    \CSI2RAW8_inst/u_control_capture/wc[15] ,
    \CSI2RAW8_inst/u_control_capture/wc[14] ,
    \CSI2RAW8_inst/u_control_capture/wc[13] ,
    \CSI2RAW8_inst/u_control_capture/wc[12] ,
    \CSI2RAW8_inst/u_control_capture/wc[11] ,
    \CSI2RAW8_inst/u_control_capture/wc[10] ,
    \CSI2RAW8_inst/u_control_capture/wc[9] ,
    \CSI2RAW8_inst/u_control_capture/wc[8] ,
    \CSI2RAW8_inst/u_control_capture/wc[7] ,
    \CSI2RAW8_inst/u_control_capture/wc[6] ,
    \CSI2RAW8_inst/u_control_capture/wc[5] ,
    \CSI2RAW8_inst/u_control_capture/wc[4] ,
    \CSI2RAW8_inst/u_control_capture/wc[3] ,
    \CSI2RAW8_inst/u_control_capture/wc[2] ,
    \CSI2RAW8_inst/u_control_capture/wc[1] ,
    \CSI2RAW8_inst/sclk_l ,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input \CSI2RAW8_inst/burst_done ;
input \CSI2RAW8_inst/hs_en ;
input \CSI2RAW8_inst/term_en ;
input \CSI2RAW8_inst/lv_8bit ;
input \CSI2RAW8_inst/data[15] ;
input \CSI2RAW8_inst/data[14] ;
input \CSI2RAW8_inst/data[13] ;
input \CSI2RAW8_inst/data[12] ;
input \CSI2RAW8_inst/data[11] ;
input \CSI2RAW8_inst/data[10] ;
input \CSI2RAW8_inst/data[9] ;
input \CSI2RAW8_inst/data[8] ;
input \CSI2RAW8_inst/data[7] ;
input \CSI2RAW8_inst/data[6] ;
input \CSI2RAW8_inst/data[5] ;
input \CSI2RAW8_inst/data[4] ;
input \CSI2RAW8_inst/data[3] ;
input \CSI2RAW8_inst/data[2] ;
input \CSI2RAW8_inst/data[1] ;
input \CSI2RAW8_inst/data[0] ;
input \CSI2RAW8_inst/u_control_capture/cnt[15] ;
input \CSI2RAW8_inst/u_control_capture/cnt[14] ;
input \CSI2RAW8_inst/u_control_capture/cnt[13] ;
input \CSI2RAW8_inst/u_control_capture/cnt[12] ;
input \CSI2RAW8_inst/u_control_capture/cnt[11] ;
input \CSI2RAW8_inst/u_control_capture/cnt[10] ;
input \CSI2RAW8_inst/u_control_capture/cnt[9] ;
input \CSI2RAW8_inst/u_control_capture/cnt[8] ;
input \CSI2RAW8_inst/u_control_capture/cnt[7] ;
input \CSI2RAW8_inst/u_control_capture/cnt[6] ;
input \CSI2RAW8_inst/u_control_capture/cnt[5] ;
input \CSI2RAW8_inst/u_control_capture/cnt[4] ;
input \CSI2RAW8_inst/u_control_capture/cnt[3] ;
input \CSI2RAW8_inst/u_control_capture/cnt[2] ;
input \CSI2RAW8_inst/u_control_capture/cnt[1] ;
input \CSI2RAW8_inst/u_control_capture/cnt[0] ;
input \CSI2RAW8_inst/u_control_capture/wc[15] ;
input \CSI2RAW8_inst/u_control_capture/wc[14] ;
input \CSI2RAW8_inst/u_control_capture/wc[13] ;
input \CSI2RAW8_inst/u_control_capture/wc[12] ;
input \CSI2RAW8_inst/u_control_capture/wc[11] ;
input \CSI2RAW8_inst/u_control_capture/wc[10] ;
input \CSI2RAW8_inst/u_control_capture/wc[9] ;
input \CSI2RAW8_inst/u_control_capture/wc[8] ;
input \CSI2RAW8_inst/u_control_capture/wc[7] ;
input \CSI2RAW8_inst/u_control_capture/wc[6] ;
input \CSI2RAW8_inst/u_control_capture/wc[5] ;
input \CSI2RAW8_inst/u_control_capture/wc[4] ;
input \CSI2RAW8_inst/u_control_capture/wc[3] ;
input \CSI2RAW8_inst/u_control_capture/wc[2] ;
input \CSI2RAW8_inst/u_control_capture/wc[1] ;
input \CSI2RAW8_inst/sclk_l ;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire \CSI2RAW8_inst/burst_done ;
wire \CSI2RAW8_inst/hs_en ;
wire \CSI2RAW8_inst/term_en ;
wire \CSI2RAW8_inst/lv_8bit ;
wire \CSI2RAW8_inst/data[15] ;
wire \CSI2RAW8_inst/data[14] ;
wire \CSI2RAW8_inst/data[13] ;
wire \CSI2RAW8_inst/data[12] ;
wire \CSI2RAW8_inst/data[11] ;
wire \CSI2RAW8_inst/data[10] ;
wire \CSI2RAW8_inst/data[9] ;
wire \CSI2RAW8_inst/data[8] ;
wire \CSI2RAW8_inst/data[7] ;
wire \CSI2RAW8_inst/data[6] ;
wire \CSI2RAW8_inst/data[5] ;
wire \CSI2RAW8_inst/data[4] ;
wire \CSI2RAW8_inst/data[3] ;
wire \CSI2RAW8_inst/data[2] ;
wire \CSI2RAW8_inst/data[1] ;
wire \CSI2RAW8_inst/data[0] ;
wire \CSI2RAW8_inst/u_control_capture/cnt[15] ;
wire \CSI2RAW8_inst/u_control_capture/cnt[14] ;
wire \CSI2RAW8_inst/u_control_capture/cnt[13] ;
wire \CSI2RAW8_inst/u_control_capture/cnt[12] ;
wire \CSI2RAW8_inst/u_control_capture/cnt[11] ;
wire \CSI2RAW8_inst/u_control_capture/cnt[10] ;
wire \CSI2RAW8_inst/u_control_capture/cnt[9] ;
wire \CSI2RAW8_inst/u_control_capture/cnt[8] ;
wire \CSI2RAW8_inst/u_control_capture/cnt[7] ;
wire \CSI2RAW8_inst/u_control_capture/cnt[6] ;
wire \CSI2RAW8_inst/u_control_capture/cnt[5] ;
wire \CSI2RAW8_inst/u_control_capture/cnt[4] ;
wire \CSI2RAW8_inst/u_control_capture/cnt[3] ;
wire \CSI2RAW8_inst/u_control_capture/cnt[2] ;
wire \CSI2RAW8_inst/u_control_capture/cnt[1] ;
wire \CSI2RAW8_inst/u_control_capture/cnt[0] ;
wire \CSI2RAW8_inst/u_control_capture/wc[15] ;
wire \CSI2RAW8_inst/u_control_capture/wc[14] ;
wire \CSI2RAW8_inst/u_control_capture/wc[13] ;
wire \CSI2RAW8_inst/u_control_capture/wc[12] ;
wire \CSI2RAW8_inst/u_control_capture/wc[11] ;
wire \CSI2RAW8_inst/u_control_capture/wc[10] ;
wire \CSI2RAW8_inst/u_control_capture/wc[9] ;
wire \CSI2RAW8_inst/u_control_capture/wc[8] ;
wire \CSI2RAW8_inst/u_control_capture/wc[7] ;
wire \CSI2RAW8_inst/u_control_capture/wc[6] ;
wire \CSI2RAW8_inst/u_control_capture/wc[5] ;
wire \CSI2RAW8_inst/u_control_capture/wc[4] ;
wire \CSI2RAW8_inst/u_control_capture/wc[3] ;
wire \CSI2RAW8_inst/u_control_capture/wc[2] ;
wire \CSI2RAW8_inst/u_control_capture/wc[1] ;
wire \CSI2RAW8_inst/sclk_l ;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;
wire tdo_er2;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(tdo_er2)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top_0  u_la0_top(
    .control(control0[9:0]),
    .trig0_i({\CSI2RAW8_inst/data[15] ,\CSI2RAW8_inst/data[14] ,\CSI2RAW8_inst/data[13] ,\CSI2RAW8_inst/data[12] ,\CSI2RAW8_inst/data[11] ,\CSI2RAW8_inst/data[10] ,\CSI2RAW8_inst/data[9] ,\CSI2RAW8_inst/data[8] ,\CSI2RAW8_inst/data[7] ,\CSI2RAW8_inst/data[6] ,\CSI2RAW8_inst/data[5] ,\CSI2RAW8_inst/data[4] ,\CSI2RAW8_inst/data[3] ,\CSI2RAW8_inst/data[2] ,\CSI2RAW8_inst/data[1] ,\CSI2RAW8_inst/data[0] }),
    .data_i({\CSI2RAW8_inst/burst_done ,\CSI2RAW8_inst/hs_en ,\CSI2RAW8_inst/term_en ,\CSI2RAW8_inst/lv_8bit ,\CSI2RAW8_inst/data[15] ,\CSI2RAW8_inst/data[14] ,\CSI2RAW8_inst/data[13] ,\CSI2RAW8_inst/data[12] ,\CSI2RAW8_inst/data[11] ,\CSI2RAW8_inst/data[10] ,\CSI2RAW8_inst/data[9] ,\CSI2RAW8_inst/data[8] ,\CSI2RAW8_inst/data[7] ,\CSI2RAW8_inst/data[6] ,\CSI2RAW8_inst/data[5] ,\CSI2RAW8_inst/data[4] ,\CSI2RAW8_inst/data[3] ,\CSI2RAW8_inst/data[2] ,\CSI2RAW8_inst/data[1] ,\CSI2RAW8_inst/data[0] ,\CSI2RAW8_inst/u_control_capture/cnt[15] ,\CSI2RAW8_inst/u_control_capture/cnt[14] ,\CSI2RAW8_inst/u_control_capture/cnt[13] ,\CSI2RAW8_inst/u_control_capture/cnt[12] ,\CSI2RAW8_inst/u_control_capture/cnt[11] ,\CSI2RAW8_inst/u_control_capture/cnt[10] ,\CSI2RAW8_inst/u_control_capture/cnt[9] ,\CSI2RAW8_inst/u_control_capture/cnt[8] ,\CSI2RAW8_inst/u_control_capture/cnt[7] ,\CSI2RAW8_inst/u_control_capture/cnt[6] ,\CSI2RAW8_inst/u_control_capture/cnt[5] ,\CSI2RAW8_inst/u_control_capture/cnt[4] ,\CSI2RAW8_inst/u_control_capture/cnt[3] ,\CSI2RAW8_inst/u_control_capture/cnt[2] ,\CSI2RAW8_inst/u_control_capture/cnt[1] ,\CSI2RAW8_inst/u_control_capture/cnt[0] ,\CSI2RAW8_inst/u_control_capture/wc[15] ,\CSI2RAW8_inst/u_control_capture/wc[14] ,\CSI2RAW8_inst/u_control_capture/wc[13] ,\CSI2RAW8_inst/u_control_capture/wc[12] ,\CSI2RAW8_inst/u_control_capture/wc[11] ,\CSI2RAW8_inst/u_control_capture/wc[10] ,\CSI2RAW8_inst/u_control_capture/wc[9] ,\CSI2RAW8_inst/u_control_capture/wc[8] ,\CSI2RAW8_inst/u_control_capture/wc[7] ,\CSI2RAW8_inst/u_control_capture/wc[6] ,\CSI2RAW8_inst/u_control_capture/wc[5] ,\CSI2RAW8_inst/u_control_capture/wc[4] ,\CSI2RAW8_inst/u_control_capture/wc[3] ,\CSI2RAW8_inst/u_control_capture/wc[2] ,\CSI2RAW8_inst/u_control_capture/wc[1] }),
    .clk_i(\CSI2RAW8_inst/sclk_l )
);

endmodule
//
// Written by Synplify Pro 
// Product Version "P-2019.09G-Beta2"
// Program "Synplify Pro", Mapper "mapgw, Build 1521R"
// Wed Mar 11 15:29:00 2020
//
// Source file index table:
// Object locations will have the form <file>:<line>
// file 0 "\d:\gowin\gowin_v1.9.3.01beta_37928_20200110\synplifypro\lib\generic\gw2a.v "
// file 1 "\d:\gowin\gowin_v1.9.3.01beta_37928_20200110\synplifypro\lib\vlog\hypermods.v "
// file 2 "\d:\gowin\gowin_v1.9.3.01beta_37928_20200110\synplifypro\lib\vlog\umr_capim.v "
// file 3 "\d:\gowin\gowin_v1.9.3.01beta_37928_20200110\synplifypro\lib\vlog\scemi_objects.v "
// file 4 "\d:\gowin\gowin_v1.9.3.01beta_37928_20200110\synplifypro\lib\vlog\scemi_pipes.svh "
// file 5 "\d:\proj\dk_video_csi\temp\gao\ao_control\gw_con_parameter.v "
// file 6 "\d:\proj\dk_video_csi\temp\gao\ao_control\gw_con_top_define.v "
// file 7 "\d:\gowin\gowin_v1.9.3.01beta_37928_20200110\ide\data\ipcores\gao\gw_con\gw_con_top.v "
// file 8 "\d:\gowin\gowin_v1.9.3.01beta_37928_20200110\synplifypro\lib\nlconst.dat "

`timescale 100 ps/100 ps
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
nGQjNTRggZWOT6sWc6oyraDUFLfWAO/HbLF6wXbCqXPNp9WCDJpv1rHVczOIVgncR/b0+UeSwebZ
OxlPzCeuO1qPl8FPTKiUyycPd+J0aSTr5vl+//g43DlAnrAZWpp+9NwkyX7Tl4KQV38q+/ZFnqAd
fKrxDpwkhDu4v9GmdKTtVryneeZJtk+qfqQLeux8ui4DI7WokBCiLCcnunBZc7zPDJ4RNHhhj/d6
kphLiA+2e7BZhQi3+S17OFvZZeAZqB9QHyWn8tsgCw/p96pTPtatJ/h1TGMYgxgbBmCeWweLMmye
bCwg5pbhghYptD2zVIQFJWuiylXMfypQ3ZpFdA==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
x5gHfLwQ9h6IkqXYFQsKYOoMTbgAOviKZwc0Vf339pYT772gCzJCT3UDF+YsUsYbK+Pq7BKRT6Uf
HBulNYuf7y+Ku9k8h5gb4vT0dUa4DG8OSdHb7R0AC/h0AeBTlns2hBJ4OSQGxyyNBp2s9HonSdOM
8ZWZFAphVVtPxikUpfU8q9qzyHTb9jMLF3VfqHt1hy3qcsmu5t+UPmv9c2zjTl4NXRMUl5483dXo
fMq4baFS/ju/wiHFuRhteazMg0mM6BfGhtM2aDlFaVzlnFbwItgar6Mu4Fk1u80ynR+wqXfj4ur2
96zU62Pm3UBbG8dYUGOAgfAhYDkhAs6USGbytQ==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=7104)
`pragma protect data_block
S64wz9lq30aLaC+kL/X10osfDUSymmrQf6hdQCYuLnmlW6w0Fzin4aO0g/WUobnGsoCOY7+vwaK7
shINCGen4o92p7HrSWBdN+5Baowett5dwKHQqJmKXDf8kRu2EUM6L5usvI7gmjwb0Oqr0AOxGdMA
IEt240OIHMHC5+4DWcK1R5uW4oisAZTZ0NJomTQDaMYTf0vbCXRvBfHpZ4l5DtYYykQ+1wrCdaX8
sSH+7Kja8QmLHvKxnpa8f5JIgVG/ucAiaLjJCwWMxb9Jgg651lo4it+/5Tpuo5y2qsnz4H1JMNUn
Uj2Wb4mlOEYAAuxfOQgISpA8CPBcEc7sbHGRaiqACMoKpmzuzNxNUD8P5cv6ovUqQfJUioqy8RZU
ncsdMPHyh5mNATv+rgnC5o/KV93EFFByE293XvqXEYEjt9+B0tjML3MngPfTex/cJ2bRYI1Y29hm
XTL62PjJKbMzmK9NpFeIkHzsZDbc2u2z/BIavl6tVtDLm+SAcnppavWyK/5wQreqZ2yB53u9z2o8
LprLjQ9sr4VB4syjJwQmDoIF3R2IbM/QcfbvefBq4dq5wIAzfUOIsG7ArZLpKq5bpD2Zb8A9OHiX
uvKXXGCAt2zRRcVLod4NupUa6X2EHnU26zdjJmoMtd40HPn4cS1oNYsj8oDgnMRuf/Usf2EPCPzZ
zBwI1jWvbx/LDqAKeiJy5p6Z3ppYHfexLl4KVFJwvZN/UAIWIEdE4gMnasijR0V/X7zNIff2Z+mg
Vst3itLdrWLhIpU72gmh+FTfXmgP5G0QzeUXu+8N1eSeRol7/A0ii/TmT6olTEgp5qz99PEILD9D
dwbTqx6rbR/vbvZYn5A6MKVaJHf1Cf2AGsVHwSde1kyO3hEKtQ4r9nRWUIdDLZuN0jDbKAOGjSOj
cKQrNjYtn3fCdAE+vAydqBHJo0aNdCmOVR4Q2pRU6nYrm/btQlG2q7hLFtC/KPp2DUkDmxN8r+5B
jtXBUi4kv0tFiBkb0PSxuTRWBbmxgMHvu2TByRH6BUq6yGS45JSdbjpP0iYwguTga9uQlQJseJvN
j15bPLNnu23qzXFj4YABLhVMn3u2NXCFJtuYMqFQMW1J4orX1gR/oDz9x64hSD6+sdyOMqp9gEDe
0WZRRJAd6GzrepdeVLDl8wkUL5q2LruU+iqjEWV6S9w6E/+nxR01/BtxYLYurB06WOIux2dQ288m
+GGE3sZDqGx+4Z8RhX1zXr+jWRREuhScq0o8HakXzrQJ5d6LY3XsmvevNbnVF62XHGOq0jtREcXU
H1rGoR5lC3ijAvpx7b8Nk6N9VmI+ia0y17PcS32wivatHlatOvDz21513YSpkq/Yw2A6uJRl8KVH
Jj+kLgnAtJuMsFxxnHHDEd0DwbhpHYNlklIcez4hcNHHcW8UY+129G8pPPfxT0aJwrvc8xdF3FO5
zGC7rZuAhq3x1cJ/zlTFsepDtjwvqoqUCODzgXBkdDzWftJn68ittbbm+zbQzXZHy39+5j/0bQGq
xrYRoc7uHFk9KdSbpbDJdvad2clSy0ty9w4csPYjbsz+kkb94vouUIdy2WpnMkdbST/cPwsGLpfj
udJD5z0gsk2qDLqeePnl3U/C9moYz+Cw5pa2tiYU0V8BmX7+oShtCNHaGx/694KY617H2GQzy3oA
m7axRdZFb0Wf5dz0Nx2TmDvYGlw8284EwrgIzrOmqP0aBAPXESpUujnN+olGWShGRd5EtgOyQLgI
HhCppZtOjMPSKULg1NinMUMFPFZIn3dNlRGv2wFaiFFWDgFJnKxRNHujBhtdwAf3yifrXHjvjlq+
rdBW/36IfXTsD2Hk9yW8sCyFEJ8thBI9kX8v9IynnWfRY77pExP+MXu6n1mMsAGI5+NMIIvtD3/I
8xOHQ4Fm3nw61qa/ENEbZE2xLwnNBdbKhRkOJ5E61hofSr+tdUO7JXbd6HEDKhyQgNHJRVAlCaZg
nxVNBSyNe05LUxwkXsArTwvBn8XteTvnwreP7Rvd46oUPX9at5gkj45CfbJkoid5ejxoP7oRA8pc
b+LtAJCrMLquvMjrcRKEjqw+yyUwIcTu2KqmtaORXZbFfDMTQidCAL5iiZiQBMmtRO3/2JWSeO/z
yisWQmRAJxgLaoyfQTxLqqv183VR0dQI10GRQNDUNkuSEADQyOOj93ejJfRl7bMQft7oV6nVSCuQ
y4cjRGk4zWKW0i3x9RhGpv3MBr3PSrgrf0dmtM+SQAyshs8XMHzJevWf/0Y+78vbIDJJg1KwCgc5
uDOLVwDKf4yKpJU7loF9aKfWzRojoC/RpzyT9A68n5qc+QDWvPhUBWhrKN8weI5h0z8dGcwY+9z9
yED1Ockg4xGHaqcWGGWbPa5C1rZUCPgFkHsmyLX8W66yGl24nohnk0O/GNwCNhNzhVwQwtkawho2
o4AiWfYhdFKXouZ/racJoqYuoAV/t9cIMNZEG2q8vvHIXNf6/NB3QDyyNrxBmJYSwEABPH7rCvDI
rDzMLY7dGRZ1CgyuP2Ge2RY28vqO1sN05e4EbXxxz2GQTnvAf62+oTQg4B3cMKNkFUzO4xLyV4M4
A3r8mmGj/Kw5MHLbs8dl44f+P9vU/+N7IiQWRgPdfhrNIPYmrRRw0o3UEl5GQMa7ersm2H20+i3Y
FLw9medsYw903pVmzIBH2R1YUdNrYOquqVdI3cEjOHbVLruEmC9CEP6s8mRyi9ixwNK1ZGF7StYb
lYUvkpMh/FbEOutMh2dAYwuCQaKcUtQmP3d/SMDOgrDKXiJKqE6tzq7W5TDy5HWT/Y43/TdUF8BK
0jJX/krAu+lIqq+KfAkrBVy1aZR7TVrpuJptvSWUogS/ZKOQecBI+DScbiM3p7ZHod5X9Hlt+on0
Eix/WyX6Xh7Qr5AqZcNwvF6rTmcIBKjZv6j+y2Flnb7VMqDsTB8bAOoBRPnWW7yEWyy4GXrxoX8F
Pj4hlK/sGSmfTI1ioE/HOfBGFUrMTCaxpq3uOcMxBQeeNoZJzL1HfxDFntp0z1s/Rv/KJcGluUaU
LRAaH/I5r9XgOinwSRcjpBrxjS+uiwZXJu1JuCQz+pQcsbsP1hc1ZM12XHKr/G9/xkPgzCiMVkLk
E0wlaFyCxuwgxb889oZCDYq+huWYcNbgMGyi0aW+QYuE8Ha9YlNJf3A3XJxk8tTaxhWqXNp4THVn
ZU7UM9mZwAvK6ef4+/UugG5R0gLQMPPSa4+TeXQDgSYeCOWKs8fwhKrEpzgFgoPv1e20fd7MS/bU
Op1AIbsXYQcxcPvkx9+QPszLjD2V5z1vmt91ndI0sgzflNwbUVdkhMwrBYowMnJKdCru7q6mqi/a
mCV3l5rBjDVHh0LiICc4jMrrSo6EiLhNwWFJWowZWTCkUNIZNUKegYjpBs7gmpuwndeGNxVfXCZn
iVlTRNTIfWj2fb8GIQ/mJDa7hzFxv/21KhESvnTDuaEjy9HaxR0+OljsYi6owDKtW/cj4ei5Khnn
kKXigqdMoPQnBBy5+Dlu8xs2AWSIQa1wUyoGqjBATErO6LXslghIbgq3y3ExZTY5kf7IKKLBmQaz
YxJh3X/LJLQkgk7ePJveOrVRNEA1BMm4TdqAFj4pBlAUeMcilNPhQ+gX38QGT480Pc2RFSWW1+ZN
oefjAnTTwBcZ8z5Yac/0qMttIH0mDph96GRuSx8VEpQ0hr5VAkTVoUohABBRUHcb9Ls90mRafwUA
lbI3mwbhRsCkcsDJB4jutp3wOCt0BVnc3b2+PBN7AjQRSASl93ofLhAxfVQ03l1nSibvSWe1+wbG
2dUJy5u2M55OD1N5tEIcI6o95cLbNOx36bQSpDSigg8keHtqgKYe+fFnQZUWWXohOI5mATn5hRPV
KiZfXbB31Oa5A3DDm+jb5C4+D6mSI2LLcQZe6yknElDChlD9GQhlBTqUAG8cGVwlMftOZ5E8BwPe
rkBZP4Ih+w5WxPnkeYmydhqWLnoSSI6HIFK+gkJzsuTlBOU93wYBBG6Umg67l3bAjI4Xib3N5jiB
ZbFxokxItCnNtf1FFaLK0+2KHPTAPbuhOE2o2IYQpnab8Zegs05TYPyRSf2/7WpTtkDdiF7ejKlc
sPA+xM8N6R6Yrwakae3dS+Mu2Y6OntbT4U51BJmslkUEf0mWTY96RF1BVKUL5SVRgCqHRAeMyHaz
qHvSApD1czKbgf4i6g3q68umeUXAJJLiegmNd+yLjbdIGrlofjvBhlw3n6umwbU2Sqxw0NQM8HQ5
K6XxvdnDQ1OBfko4XHIFhhkhse8agYli7HJ0cpOsC0vaeHoA+BTC0lAKOkOLLD9Q+wI5y2lOBRUI
R/+2kC8ndhlEWoROS1M+bMQ8AURisonhvfmHAt62wu6CSGlbYwkp1I3sUxtx9kMmPnGSe5NHe1Jr
wGSchJ1g/D0weviUf/8UAtojoJiQUi/eezHzww2DQfz5PvREUkVQC1Se72W8wF2L4ATqFFaua12b
wGFTzC1JLsaMMaPmL8v5S0d4vhhorHtY4uzrMjEeS8uzcjyssxaVOE/ZLklT7bX8DKdlmIhWRAKV
qHHvdKv7weZ9yTsxXKWZaUpg4MHP0v0gdGecJ8xkSageBrXGZp1pI47y6W0v7bc3EMyt7rV7D2nM
hwUGuqQhktdwoQiLapiHCtuLi1cKGeScbabmqW0gFXV5ooMTafetu2mHFAhx6q02YZAPQhfcosP/
gwCqIcK1YPBEyJ60SkW9/KGp/K4XCOuyqgbcI4RHUPXCHgI8cVy2pRTbCRMb2mi3xA/Z90FEU3Xj
uQrcGrPom8pyR5E+2+9LpynAldtSRq8Zcv5RDP9JX5UzC46Wz96g6N+mgtkn2HEf65hkGMeE4lHl
7QkSgTEPQU95gFeFdkSbRIzkbBuFoYeLSRg+C2NVZafssUKr+hmVdhlxpaBI8H/Pm8bhBdMuTDXe
baF4PjmAlt+jvXOW//65RpWxZIA7UMjfPM0qvzyqNa1pxutYSAlv2o1PcmRbP4FWJgREZrqHDODh
tH6WmdjzAX/aekH+OByWGjNbusM18D6S4LlsGX3TIzolLYTrISa2x6rD/dhMH42XZ3f4Euhx3p81
JBGaLYR0T6RDiPaxX6lS3M5S/iCG33e7TN4pN6sgdSsnC1dGZG+R0hxlKTJ8/uV4NNtzkPA/n3Zb
V/Ygx3XbsyC5jh+IHQvpMLdvbbZi3eiwvHwY5FHbhbBG5/UA8B1WTNIozV+Inb6mH6Ql6upBbU7n
1BfBMCH3b7kgLpqj8FycR6TbdsifLKegykv4rvvIUfrFos4NRkDaZigtCaiIZnVXVpTO1pWb4zif
EgNlCkNstuHrqcoEPD3crhgsmeH6Xf/rz8L/q1j9Kgqpq9qPUwUmttjr3ADtq4sTp8OgyDp2JaY4
6vYD3iIlvsrZsntzpWMm6c9TPsd5cTVpBnUWd7aB7v0eMN8BEbrJcwZPQef53ogY0XqPYaEL+gko
csex+bKwfWUBCIa0CQFsVSMTJe9XfCiItiSDI5COuXus8rISVFLgwl9d8kiYz0wW4Uc5/jGhwGVX
zhQTdRp0cN9HA57fWmind5vjXwI0qe9yRK78v1upOq1Vmms4KMz/teObjCkPbX2B9HaUQiRhVt33
tNliZfjsVNVTY/oHA5nCz++NA1vN4U0qKQhI2MagqKVuWvCmdyqLP+lf8FTnYwrGXYeg4MOZ0T0T
WzhUhv2C/dNmk8N6/bBUkJuH+WXhb1pveUkLBM3M3YQIYKbjMZTNooiG8dvzTIWbZRipW0rfltGg
rxX98Xl4nw43GXLStEFK8zFBjSoYFqVRMrxgyT+1VKGR8kEYIam3L1ZeP2qWvw7+Yv6+8rFZzKeZ
fVjENVwZ+10eIBH9pHtOZtC8NMv9St1efR33q84L3UZ9YoN+brKClkspTGiw7xM6WMZxur4Xj5K7
3Ct95Si7wTDo7hrfsHA7EZhyCAu3CDJg30Yc8iHhD6oCXL5Jbn4cgi0JAiiIUmXu0lXra4o1OrJG
OEmhCcpHIaRtlsDuyhat8zQI33wGe7LmOThpLb65qT3WWK5DJVxnJb+BNALWwz0bNckMVcWjPjvZ
wbWRKCo3RJNQXFiYWGpDlujc/LoTckBnG42+9RtV5FteQdb3k2KWxs+EyDzmWuwJzt9tmff0eZZC
gktiPz3lhmWywZtI/GZY4E7D6zOo8f/Gou79Sll1LmKjrJoYerB7+BHDEkWr6bl+uR6LvuCO1NMh
8G/+IcsgDLbpZB5T0XfebVnp9EkfVSklT21oxBixgi3KSFOi9eWAJp3zXrTY4RlxpBXcMTr3gvlF
chOj9VsyNQAX9jp8eIZrx8UAZf0uBe5I9WVQ0cOGJDdwumtgdvmAwYyiHwzyGNZ0lUMkzKNMQtXA
2Gf0xVP0mkRcezCmiqoFTGu35veszVCnM+LYQe9Vf18LaD4Cv2ztI1+RjTTn996RNBHkUR0n1ZVR
/JOkPTQGZ2I7wRc+UDlZlZgbyPSSfBJJjoDBUuNGacDYSB5RMhrmKwpu4ej7ESSqnx9xiLQRCJ8k
mhlxgHN0L4RyNYLHfuQNU12gepUGGjy8CgrLxeV3SRDIRuWqMADgfDgLrypwBqPorM2sMs9ptX68
ktZFXcwxJdcqo7diINqZGmGrlEIfuh4cTGp2j0BMfMgzbeYUpfaMOC90U66LKoub+dp7aaBdyyzX
OSl858zl6Lw6wD+bMtiqGboc18KwIF7NyesiOte1SF1CjCbIawvMNlAO7ORmQ5RZyOUKgnkOiTBO
3vgakwZXogeXnYrZXjwAKHlPuWAmiiXRs1sBu+slXY6MDMQv5sp6AAd4wj5DD47Ekvqa49Im77Pl
NnCFOod0mtE0+999pgisGX3rlFq1CqsapTgnX4XvsCrYQmxZsdAdIbjiQxIWZZGwy6zAFPi/YY5+
l9MTHXZBO8G1+iJtEENsF/RXb2fdkDj/p/VhmljDFL5DsGk7Iuk+X8OrazniOoDPqXtFaPPSb8d7
o5CwXbtQMmuthC+kjoomZmrJ7SmFneiw9p39ckPoZA2RqgYsWYTMD0wcwAsTHe8T32VGjAxHXb4w
vTIAVNH5wpxDKNOAodjFMSwz3qBcghDJwctosIPna1U3oU6paurBSDH1fPESGHShTsuCDPkNt/3A
ymgFnsOCYBzu6zuo/jECemOIMVLykEINTED/91fxnmmgmX0J0flYvVtq4MNZ7qWX/Wo5ssrMIMkz
+US0P2+t56X9yc9EsClGzRzNJdSAzFM6c2jZIz+p/VjrgKuyT0lhQPWEw9G2WUpB4xTtPhTsjQ6v
mG8o48RabcM9zOjLqYSQR87B9BHH2pD9pf5QtXTDjkGO/b6++aycn4oNCN+v+vrgGJAEHC2N13cW
RRh+i/1eIU5DUwBhFf5WegUCuhV5e1aNoLzmgAGOTf1evg5y7IJfTgg0FsnHXgMwBEYgCtiAEjLe
0+Fs1Yd0yMMl4q3DKH7wVIpZQBeYYVM+ENr8w9U8jS8N6q0JPGSbCNA3GQaqtZvsL4+RiJrXe3xr
vUIoMnxkHHR+ix3y/23R8hvVvhnvOnx/0YIB0fBy/ema0AnH+iBSjFaYLM7vuJvyCr4Q769jzT5q
u7RGBNQo8mXXoFmEe/suMcTSbeSuK/hwYB12bAyIDoaLToVOhHryyR514+pQCMz5KgS66TV9D3oi
a/3e6C0Og1t4KWg6it+TGLGw8RGJPh0MXoqR7y01no2Rpjs7MzlLH3E3IYZambc9YpdbtDCasv8W
Q5wKK2d9xr7MAU9XOTwscE4Xv9d6cr/bfirH7Lvjg2LWz6KWEu/UAn0YQZ+V/J4VsTn/bVrk/eaX
PZpSsFSesf7JBcYVGbKbmSTCH9iYA3dW//LvyPXuTz5V3686tABQqe521AR3OcVGr/2VHkbt1upz
PvROv6o6kNCj7NZTUGGkn4ZIjnqqhPuDPqHlVtHGN3t0V02WlcB9gqiVB7Z2sGteiBHKp/yEXja4
WbAWTDyJ7DqA36BuJwDo3vAQFDA8/dAvepjqYD5r5VqbJqudRyjsHuOLEKbdtJGZm5zWvGYYoNw0
ARqR4aiIMMSp6nIJUdiKc0lWZuie+ubOIBGZoX6OjWbm6NGTODFAD61hWGFgoR9yL7yhLuMtcrGg
1TKst12FTuVTDpT519TrwCAavJu5jLB6vVooDxUWfZRhgJOub7NYxx2A4aj95j5s8TuFqqdLPP0T
H41qe26XL2EUnRsQDXFX/JkHH/mNpXkNxNqJz/c7h08UTGn0tsEMypIkGYBirhZWkRC6YBrKAjzJ
NkVXRmNFKCPFwh7DsIYwq0hUjS6fd5KB4Sh0Go2a7t9nBhMVMr5R9QHyQr/CGMKLzvgpaxXTpHR0
mTkHjJNAeWzNVdYzTWG3sLqhC/9dFOfU6F3FLuN3WlsEkpyv1vPQ9iGl3MND2k5O3dPIxobPRmf3
o0T1oRw3gEQ1Kj8777jZO9I8Uny3h5KOv7pbKlOWeCjWb6MJ6N4Ct0TDBq++Skyv6YJipDIhJKqa
pL9IgvVUPM9ZtveUpCFTSnLh9WPRuJOTkQoYQkSpyPQuk0z06SOUgBU0Oasif2RC0ZOhOUlalUQ8
iWlh08Dv79eNGZIHJ2wstW67cX6d2mOR1u8UerxZXwuOWv9t/tKoUYlGruZ3JQ1LwWVlk4y2K7/E
cXY9I9YCQPJrMV7+Us2RifXM900SRft/vmFecRAQ2L1Fw9cy3hd7YRBcUpf7fL5s3i0a11xQQxXB
fKiiV+Dg9Xj3a7HX/u0bcnQ2VDgemdvOJMw2cNl/Q5S6zTYjGpvaHwFCd/46YWACiRCG/5cKoN/N
ueBzxbkXfVAkf9VJNTy85ep1a+NzjfuaU58ahtvTO9miRK2ZbucCsOeak61+6CIbB2es45bLzRml
6xUZSEsRZDN3t+uvmw/ujPADTmMzltXFpRqu1MmSaudaOK2aDXAZJj4/t1SdaNwAi4rMr64MWCvM
8GSpZVXHAaQ9MRoomQALFHzCNXBftQALac4Vm154Rr9JdfpO+C2zRAS2zrv0jBukrxc+kjOwKyJ7
oAKfYroPTvkgcIknimdNFqohPzHvcSroA3qsC5aJ7jnQEYtqbko+0p+U6cC1i/x7G72SPOr2cWep
jMkU1vNJv7a30OSBx4zak5x6FN78jTeGb4CUaxVMBVHzpYdqllvYP+7PDZeZ8IJcJb9VHzWWL+Vy
SvQBtEM4uwrUSG6Bo8Ecj3HBEktuN33NYSeSPXzzuMySZdAALD6Es2xXigIVqPCQceUDCVOe3BlK
WHF5B9WHHOL1SmhGO2VBaGYunZCbeQdtI5p0jnTVH8yXQHq4WzNk/v+igL4NWTOOs4Mp/prj+wkE
BCttwh96l3EqP2y27GcHnn6z4FYKMueLuhDDh4vSVAReMFkyObjkr958tFwKukAg05mM3Pgh/LmX
3PzsF4PQXOQizNvIyNLkHZ3B6iWi8rtPs4KQKEu5ZOsbQC+9
`pragma protect end_protected
//
// Written by Synplify Pro 
// Product Version "P-2019.09G-Beta2"
// Program "Synplify Pro", Mapper "mapgw, Build 1521R"
// Wed Mar 11 15:29:17 2020
//
// Source file index table:
// Object locations will have the form <file>:<line>
// file 0 "\d:\gowin\gowin_v1.9.3.01beta_37928_20200110\synplifypro\lib\generic\gw2a.v "
// file 1 "\d:\gowin\gowin_v1.9.3.01beta_37928_20200110\synplifypro\lib\vlog\hypermods.v "
// file 2 "\d:\gowin\gowin_v1.9.3.01beta_37928_20200110\synplifypro\lib\vlog\umr_capim.v "
// file 3 "\d:\gowin\gowin_v1.9.3.01beta_37928_20200110\synplifypro\lib\vlog\scemi_objects.v "
// file 4 "\d:\gowin\gowin_v1.9.3.01beta_37928_20200110\synplifypro\lib\vlog\scemi_pipes.svh "
// file 5 "\d:\proj\dk_video_csi\temp\gao\ao_0\gw_ao_parameter.v "
// file 6 "\d:\proj\dk_video_csi\temp\gao\ao_0\gw_ao_top_define.v "
// file 7 "\d:\proj\dk_video_csi\temp\gao\ao_0\gw_ao_expression.v "
// file 8 "\d:\gowin\gowin_v1.9.3.01beta_37928_20200110\ide\data\ipcores\gao\gw_ao_0\gw_ao_crc32.v "
// file 9 "\d:\gowin\gowin_v1.9.3.01beta_37928_20200110\ide\data\ipcores\gao\gw_ao_0\gw_ao_define.v "
// file 10 "\d:\gowin\gowin_v1.9.3.01beta_37928_20200110\ide\data\ipcores\gao\gw_ao_0\gw_ao_match.v "
// file 11 "\d:\gowin\gowin_v1.9.3.01beta_37928_20200110\ide\data\ipcores\gao\gw_ao_0\gw_ao_mem_ctrl.v "
// file 12 "\d:\gowin\gowin_v1.9.3.01beta_37928_20200110\ide\data\ipcores\gao\gw_ao_0\gw_ao_top.v "
// file 13 "\d:\gowin\gowin_v1.9.3.01beta_37928_20200110\synplifypro\lib\nlconst.dat "

`timescale 100 ps/100 ps
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
DI4rXVSqQQakdxUiFbNMpUcFqLtxiH/v9VC2fotO6RT5oJx4ujfd+d8ntglwi9SznfUhuCDdANfH
XYMgV7tqilOQ2ZawjyjFzCrZ5SPXrGgsruT0nRljnPbi6qkiFtugOcQTRLawx9T7//cBM+KloXTA
NW5UEesUVY6XIevfIUZGJ1ure5Ny3juAG8DwrfgVKoVsVbpFHGqkn14/CuCrPfgd3cNIeMnz2tdU
fIIQcJuw7/y7oxsPIHnSNjduB2VlABUbTul3/U+MLlIz6QrQXnGGd0gsk0VzmjNw5t92AUKNXFJQ
KgZfLCLpjgQ/ZbGsMSNTxIFdLQdlxHMJmC0vaQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
BJq830S/kOcQBA2JJ2q4S6I8jB9jjQ+2w4M1vD4Tqw23sKPDOhifxjr0/o3W8kskkjrPH5ExmJnx
4+Ax8NsC3/y94RfnMYtaR48dVDd/uZPC+H97z8xQbMlRtAPIPBxmvbm2XF9esKwvNQk33qXslMT6
Af5S+VRtkbzP466p8XNJQwyztsU9oaM7FXV1jV3HosbJuRzcKVPEOmo4Dn/DOSxaP8rd5LPjoLqS
+itgiiOB0/sBM3oF4lMqNh90Lt7h7dN75Xc5z0AOiCtIi7ReGbnoPIxpLrTX3YY2f7/TaNJjwe2m
A2muDv33kmPJYj0Qn1mVE7WUxAUWY5au4KLJvA==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=41696)
`pragma protect data_block
3l2m8UONmp/7H9fdVZbpxpmXcLOYUQ8E9OKnRpvBGbgnt6ZUHvcId2kxEzaAxjvFxStSV4e6VEkt
46PjNGDNs3ytS/kI8YaRwlrW6igEyWlDKtRlLjugAwbDVQwt73Y7FGrSExDr+8KbyvLPKAAl7cqo
OYPw66Barh7X+JCntsjtzG1wNj1Tw0M5PcFFx3lqtyyo8w9uN/URZfs3YsnYM2lWOvnHbwdieW6R
SniTaruAhFALrQyZyUcd3nBK9T2QWAowWnLfPmtqdWmCdqSOGYAHBGn4unbSX93fVAAl4DgoCEpF
ygi9DAZcykBXvh+M/yUulrl5zKZ63cn/91FNF32u3J301WUeEP3uneO9unOEP0I3oaBC61Mz+WbG
tRRkWX7avhm+XASQL/BmPHxnJwhk6Gu7jLD80SpATZlwii0QpEOmbRJVlj18udFN5bjFGFgNCebH
UyHv73shKiAAMwacQy84PpvCT/aT5onok+qLn3zskXuQSMiC14JIqOX6KIwnwOam2828G0e8N2h7
dE9wZ6D/K0Bsm1O4eMayR5tnNYLlXAf83ad7y3FWoQWqFwfIlCTHuulWmg129EImXPgzBfryCYd8
eiuxpRnkD1uWmPEoq3GDl9m2qwnSYu64dNaMC7Ui5K2TgQP0TKbIVpAnUdwcAREsiFUukyrqIi8T
z1uXCHfBHLPWkbPLuBTa598A/QDdd1yPtBN1LMppPOApMRzWMEFwApI7Mm2wl6slyLjBHj6hgAKo
ZFTVMZrjA5SLqBxjfzkXj/4r6vdO7aH7IhplXk7w2mpkVVaE+GuGyFjoCoDLn21mlPac7FJZcU3T
S2DqGCwr67otVqfP4PGHRCCFDyBknxPGvWu8xcda+B+HDGTDH+2zOOQbA/3QFaJofnvs+OUSbR2+
Bi14goCb9NH23v/MUnEGul7rAEsWqZqvCqxAILwW62ZiirXqzqLaQiqqZDup7d8ja4YWanVDD9g0
zu8fGf/GC+xO9RuY1hHzpHSP258FVrfzJXqY1WQ89avC1OO2JAOJlQT3uvtlLxTwjCLVL1Uce9Sr
fRlAXIHGKtGYBetzHk/whEk4xV1ClFrkwQms/Ds+T5kca6tP8LYejElJcapK53OCKP1M3m/hSkpK
3EG6LPix/FnSYF2o7v2bgjLckFDKCf3TVhw0an5iE2gj5yB5WHM5vgXxMFPhoBUgSdi+kmBOP3Uf
9TwPzGtsjcXxbiKjcR6pzIRvJdnpB3QpqZweJSAdiRXptFE5R6lgQha6FlI7XllY1iopvGrUGcg5
8/xKCToYn3DfoYxbanVx0UJAgJt7GLMOd1aTZB+TQfrcFzSteZFbGQ1g6GeE8y5gH8DqzZfKo0R+
WeANCzx4VCYqTVSnTBTQYcO4ocrGP9PG2j53DGpr2V0p0/uxod0edOgAtUxj5UO1L14Y5eBbXi4W
/AOsqS/msoPWdiF5JBanVA5M6BxlDH1PKGyu+86Jyxgb0aSr/6GX9lqV2anTJDMTYgzYoM7NI6rz
2C6dMoFxMTZVlJm++Ls7dKAk6ixzj4J4Nspx7Hp7VNMUJGIPZ/LwV/yY+4WoqMdp+DI4xOyt1dns
EhwfOzlztsjjqXyyYnPpPlOdzibNiMBHJ4t4JjnmXRqfDPqQ4fJRlDH9aXzKCVgjZ/Ie5lK0NBuI
gt8Lo86kpvP8Zljoflzc7QwXKFHARUjvz/pYemQX2fNtuqhGAYrXTxuA/Or/D4FXbW4gjXyB2gJi
oAYGNpxMZW39jBOSo1+fJ2az41SEBzYMJnhSohKMcEUVqOSvTyrsubpe+1ahb/YSFX4CxIoL7QWG
3nR5hOAo3ZnHhZDvlvUpJ6ceWS4qUl8tebsPsdpb7CJqgsSBablncGTZX2Tq72toNJLzUl0rejLk
gwGA2xLVUjSmO3qD4A15pKb4+6eKB5WXhmDz8jxkebwHBtlmqm5GZg4/KwX6BuOl1WFhMdVDIvFp
0rfZ0A2Y7RL6pjd8SKolMMc2wAVUiW5kqLcqvrov5XK8N1nPWd6MXWSRNRB1XFSWQ7J53JZZhmue
bfbYMfY2AGBCHli/+2MCNsvM+c35uEl7wIBPf/kpNirebQI4evfp2x+SMgonLYStj8kZwRdyo7vL
7HwKX02h8xpxOn5g7pI4BWQb+VYiBrah3SsR5quQkrAzuS0oR1WDLotgeoKWqSaO28E2EH5VdhiU
p4ewQ1sZCwerzkDSwQAzpPwJsJkJ3uc6/ZUwYUyaVcvjAfOi9s5hxlUUhYsU+0Zd8G6nxWuZUxaS
dc43CKUPv1RQsY6uldAHYMl2RdTlcFo0p0vua/Yq7Kced+UFzrBqlJY4nPlLuPtVcHwtuz4KKWF2
7iEZEjUL1ntgv2VMVCzLM2G+5vZqPakyYzQYy0frmFTR/n4g2OdS11UhaqSrpN59f/mlyj+6GGh6
KkAkEr8FNY7F9LkABdcDHZfkSds64N6OXkzt+H8AmmIH1iRzqzqqIEHheiYa7Y/8uyb30wdbQzIN
AwLNAurEM8LXRQgSB1H4uBPpj52hhY8jkk1K/NfXvh6jt5IDXtob3Ax+7qcNcnWdQPuSB07kM+HW
Nc9rYOqldVkW6AzXFALjmKkLehm887b3LeTsdLdf6p3BFYfLZyNTqJAvQ3jjHxfydbfla3Wra8m4
Q4xaAzXE9qEEyyGY3CFl9UWIvRhqzUrmEzOn9g0vfyRaC02I2soLvuZfrgNdphbZo2hfy2O2HddQ
YwlDv0XPnay7lKD0lfAvhcb85AYlZqJOJ/g1fTPbwK+Cy4kgZy4Ars7/vXIIzBQvdZUtXPzm36vd
9YoOSNrsk5LFPYUN8JSsbVqCX9fY8arcjD0+9T7Du3ubO188XsNGlNI6qhgWzUfvO7rZQ3iNwWrT
Sov0iXwXE6aMYi/vnx7SsDidveq5q6JUoa4SeJ3DhXCtpWWQYt2bMQKTBU54L57VstEUkI0pFq/9
xYHF5oWImhyoEqgxU3zmIh50Dj5YAt7ii64atLdI9z7473HdwN8RExFurrKCrCQa/+neOQ44rmaU
MP9fWKz/VuNua516dY/fPIIN2CSX9O6+usztxeQplD5xno6QFbNH9iw/wWMtcY7A7WSPjxZmhvzl
JB+ZnOerj8vvmAqU8jW26zBzo7PCzwm+VyLylGEh0R9l9M2n5oUn3T8Ogw+zdGeLPOeltTy+oSAe
nvrXfaXgit6Dn9ixb3fafUIojx5eEPTnIvtDjzIJGX1BXW+cHa/IkY4FJbaaAoW6buvOrOsMxNNj
HzORs9vqEMst7IrilgUXy3CP0ffpl/LI+ZaS5vFmdI5Vn9pvwCViI0XCjoMsOIpbhbEdIHynicij
KshSbCMms/JymIq5neSo1adoDIkQ9UyVPP3GsgIsTxiWs27+zrfxCXfVPOgsqXIDqNFl+Ul8wFzf
88aK36DXBWwukG/fqajSnPjlxHqOoefFSyB/CoArG0Qdhxhx9EEak0t2giEMh8G0RsRrrSl1FPPn
huIHEiOdVwr82krgilPn2VQpK3HiRIYdB6/W6tFPcVpLyzcmYQzB9sDlmdw6sEU2IILhFqVbOUM0
D2Ve43Z/5OzdzTg6slblsneWqZXFyiS+ULHsZG5tcSL18mFkyZ+FDZJUpVnB1e2PtAIR7F9ZIh8M
oHYOS5iCWO15c3K6hq22Au70cbLCQxTTsURXP/6ZG2k3BIUBwHw495PCR3d2Tf/6AYJ1jahsONyP
yuS2iJoldplxI6LhNnyVwUl+gfZzSTGTuo27spBx/+PcRaYd83LuUYB4RePzki8nhAiuevC7mvx/
Hoo/JtJJjDhoghjojwL2pM9xYzSc82C0Xe5UF9o4AO2PCsDl77CSQD8oTcLc6hTX+ibCEUbhuEpy
Up+WTtLMjUa4PhBal4BTT3gxQhWVmxw2Iz8KCTW7jA/GUC6jyq8molP9Py79WpxP0uKQ55MIypaf
vCLS6upoAAZWWgXJrl5U2cgCYZqwNec20L1JDedcsRx7D6PlrXSbOhaTTYrhEUAmYpgtrXuKmsDn
ZR3w1//nt4MZUqBM/vqUluk/jna3UH3AHsKTz3nreMm/7MkrJ7d0FxrfhGPPL3pjJqmGOWBBQC/N
xFsZrAwpltYcbWlwSYP9ohWKSf7PxNFPGLYbPPSRxZ6x/1vo7Le89dxoq4wwAlhHh+IZx+UJNHbQ
0HDu70/IfDVi3y7Qu0TCXQprfyZ/sW98vXSaFOFIdLXSYp9V+aHD1bE1HnFxMfHRjwrezh7yHdEz
xDkPXVcMeQuWYBK2PpsD0mjc9ofdjAyGe1CfqIfbsa21sf7hUZYQQ7RoeT5Q9VK0rJu9YbgTDvx2
lzs1m8QBXshrOHZaZLiuI4RGW14Ig9dRzFSNfsyeL1og4KJOgO+qTNzZAslt2IKFz1PnmII+1nfQ
I1emSMSkxqy/OMoZQQC5kYhVvGk+HzQYBeR/eEnKmBA3G4PWPGvydoplgYVsMsSrLSOk+CHMPtfC
388d3PGHrVsw87mK33yRFbrXY+sfBgXiqss9/e5orAhC8iOJ3ndANTZYzp69mBETl+Q+dFp+VWR5
YaZzZVnqFAzCJWZv2kcDk1pCOSmRynYSBofB20dpGr/DsQOPYlMFm8QhNn6ceeDu6q4KFkoUcRZG
Kxye24rN/90ZluC3/9g9vwFUcbEJ5zKcQxJO8NM4jqPHn9YkOfVOMp+SPeJXrVa+TNkEBJYR/Pu1
2pN3aP7tfoTaZNKqCHgWdxPy/qRu5JQ3O+sd+A2GRjx1ruXxxZgXbl20NEk5JMW0QEBWnQD64Hpl
SM+XzJBVM6UE9Bg3NVTAGvUVlFT6jIN1TotWFbiVOoxx++Qw/Tdm3hlIiXEFpBA/cYFq/9QCdX0q
FN0tTVGHvumFN6SOBV5Pp7V5R97EivmB3ptz70v7RqW6BsrHsfqLAczCMhzBdOb8TNlCSAoJuKD6
e/Str6mk4lzD/9ENYC5zvxNd5Ruvh8Wp86cpfCNrDTDSKwxKlcSZXUARXP2miHv98avHVpRZuzw2
ZjxdKOg4FSgAa/FXstrToVuRf0rsnX9oukqfJqXxFHJf+SQESCURDMXjLpxZW3FQgt3JvvygilWf
29ltaF21wmQhiXvUnRgM+tD4gZByNQV2CYmsUCIotjNik/LspnI5YGxAKpXV69QhZkjiAAhb7t4+
0EhF2uS9/pWyegO2hEMtjlIKYCXFM1sxOXCYvEviUPRcpgnXTxQ+LkdcmUNICZYn0s9GbNvFUb0W
tfBXvZ7EGdX+LuRFELlusFn/XxtYw8BKnwNvxPDCw+QuLmxNWPZHQhuiRBa3dYHo72YLuzqPbmN0
8RUykVi+H2uFjUS5X1X4J6eKa5K/Z/ivGsXjT/tBAKCt7PvWDaRACa8Erb1qDwfchayy51md9uwT
LtoiG3l7OZdn6P393AGxVXjTRPaX9QME3cnOWdMok3SyIUqPzffStPoAC60AWesGlvDTD8m4Zf4G
7YNjtSEa5jOmfJeaQ1s3/O3bDyQmUK8DqoqJYwhQxJClqlbzsrH1137ukPprjnJEbUSVeHNYV/fO
fP2RSo7fnpmLM7tlihGQZOW6OvsLO010Y1ar/V/pYtNDGbBVeEs16b01ltwQCPX9RJBeRDzJfzKx
/W+5oHVbZm3DztY3XMhl8TPPO3ZjlhzZq1DgxoHN0faEuhxUtu5afUF5PIlUDud5+l6AYrdXfDNH
KWO4gPf00fmC7ZM7o/EtgJa3UC3a+SoDv3A75UQ1KuzIi9joMaujtKkie7fUViyw55FaG95+RIP9
IXz60suzeRqlc1TWrtFGV6KpY7LdmOLAX1CfJyQy2OUhN8WA0ruPr4x1uimzEgPQfpYAXFTgCDQi
39b97AccP5ijZgqUqImBHiLCeYcyUc81M15rfQ+FQgDm3NOJ23Z9dRMth2MMvOXo827xBl/wI1CA
Vq/+FwWg7Ww2IZOor91O/mbKPc3g+a8ewvvzJt1lhfJmtODmbHG9dS8/B91vH9ZdWsUHfW3/UNRM
0xbQuVytlk7Fo9lPsVEPq5W+2yH7Vgk/Z/88gk/15miDXi2lUTaj4ycIyYABm5yX3UJqwueHHINX
OgKuD0k2plqN+48a/JahyInwngT3X049LD6Bqp7D5bcGZmoHrMdcIcgCHcPGa6RunK0vPydTXFO0
NEFt1bVn7Ba74z+QQ67j/9C+80laJziempfqedH7YhgMNcoOTH9/IFXJuus1NmAl6AIC/TW3W4Xg
RFAw/guLPrE/J76O+0xaaEq9PwaLGdTbOZpngrOllPfCd/kPPjIsSWlzx5/ISN/4guaLFT9QkHct
gmsIfqzY/tfjyrHchV9FmcahyqbqNNLnbil3SfaGvxEwhpknCw8N/hAg19NpptobwLxR1kq1QGNh
lw2nQ5/HdEuFpjNefM8PGy7/MuFua7y2n+TUGNXxWHUt0Q3VUg71O7+yBafHDmoEFeP671f3wOge
BKNIoqNdl4GWyKsa61SqDt9x9MEkCpQFcVFR+bojs9kTILKQE5QlJCY+RoXUf9yRuWiByWTdTwkz
mNndetafLpZfnTO68cIaAdoPJiyK03hUiUzrkpo/t7oFpzPkoqmqIFJptek5eyQZe3s2zP5epXcu
ofsQPew8yVaFdLpEZFlIC74+3geMG9tws0AmQrab4Mh97ed1Z+AegyBLkhIvOtGuKLUgWVIawRMP
bLRe2dMKuQvCFZ1MsfBBmFtswXFDbyIxgQFNYU0tDI4BoO0sNBc43a+hc+MPsN1mRY2TKKbsu5cl
WdM8HPnS/d3SnxFSyxdK9eR6/gktxHBrVorKz2w/UY0vHoFOlpJZVoh0cT5K0tJj929HGx6KUys0
7cGaLhht7wOUOkFOsSqDJ4BoB7KzDPp2oNt93cvrD0gSnAuvJxXx2xtJqCKn66CuwXLkCzyNo5z1
Lq9GfJb4Uao+kAkFIFS6ZZdNx3GIUcwMVzaFkwtnRB2paMW1JfCTKq5dWzosqcdjJqupRZmwu+lB
86CpAH+qwO6y46iNF8jmzhvmHj13apQQMqjWu7WRrCv16X05SYopBEIAMrMmPc/1pdCmwzoQ+o8s
6LkTer+2rN4l8D5sf+/APmxJOdyUm0Aa3iSWScCGmVm1SeZ2rMfU/wbZ9ldH/cT6L18LoxuOPA/x
yn32dGWjXMC0390kdqcftFOA5i8NSCOGEJBs8keLTI/zs1gMELBXyC0Wera6noK2kQqRHcEhaQEc
eHikh+TqE5Igw7mjSN1Zz3xU2EPyjcOfJ2p3HfUOI9Y1T02cPlnq74xpjA+sCQXooOYY5scsabwt
kzVb+A+vK2AqMU+xdZfz2gxE/22t4zNWWcFqBAl6r6YzUd7duBic8elCVfe5sVDkuxjGwJk/9fIn
d+w2o2Udil710LBR2mMAwwkRUxJ/emwnpZVRgsspmlSccYCRotuJ8k/nLXPHP3LLoSGmGWPKwfUo
tRO7Pwhhpuwt7i2agGxVPckhhdl6gExaElfRHrr29DjCM5ekGZMC0Ywb0Bbr0D/xzMGXxjhEr/MM
uW0z01daDIYcf6FJOqRuBY1EXv4qiNMQbvU60l6+HNB8QaHcp/dXiRt4QKFZ4kXq+mL8wC4YV8Tc
UjugARgfoW8sYX/VA+7T67TCb+PqSpC2VmMUa7tkOPUjZGd3Bg3MOE4GOtsW8DKSV8HgMYRQCgwm
1nyRzVa9s8DPM2x5IVuGIU33AkG6c4omCbfykNMYInUp4UhKeMIoK7Oinm2bsuqksIfJdpZ+JwUO
Qiyzx1cdeLeU5MSyPUsaBDyxUWE+TD2EZcn4T0YvjUM3bN4ID/A9SOMgSDnOj81Th6GEyBUyplqD
WyceWpuK2+CKedCTihmPSQE6R0+e6HcaCb250B3lg8R4fcYB7f633DR40fofWmY5ZPqd4RDAo2MQ
kXpZK8+r8Bu14ZBMBYvNkbxZpzTAMxJmVzMEdDIizWNm7cXAovEKOvhmA051Jq42ELkoK4B0w347
ixzYSf5WHDyMfKTIpiMJL4xRC4dA7oGZpao5VrF/3vaSzgMflkojHqmmMpYG1BfSN9wlaFZbA8UP
FK6sEZZ6lQ4A0y8RA/JUm1vrzHsWkmMWsSlYXVlLDaBxs/1vgaK8ovgctbSX1mjyFDJ+yY97USTn
RJZ4RGfJ+kOoLZOhhYJ3w69RnQICGDox+FshHdD94SxoYdH1ZUUThDEtkJDWJxTNMiu1gWM/qf/G
N2O3H4dPI3k9dkFyreN7b0VY4RJStp6plrZnSvsMcWKbpqUVtEB5TJlnWLJW35NwMOtJ57NDLRkH
hG0p+4E/oc28xkOirBdRlUYJW4wp7an7S5PQp3pZfTy6B6RomDcjEaG/QT6w36+IAyGyAEWpj0p3
bWPjX/QHkwmL1HdZ/7gC5mxKgMl+xqQtsRr64lfRer8HK/7H/QaVO/DIlK/QuEXZ3rYKw6jHgITu
ExTADOeFRej7KK41TiCFBWZrTRIBcorcmjtR4HnS1e/AUq/JhWpwDpQcWOu2fvjkpMCuKpQ87cOW
gprysnJBXKr/mZb4up9l/+Y8dE/jdFeWiT8I2JNbCkxfJ41siYOfU1nEI5fALGwq4zLsv4FJUoiC
hkbZ1OgbnQYTo28CXh38umi+zcgYxZE5m335afXI0zNkqxrm+dnQN+WfDBHyd9Lv3tLk/dbAvQFY
0r9MbtvQHni20YHIS9oydd8ZZyuErWcFd1HCEhfDCijC83FnF8sjoe4Adky0d4ST7JmH/EqjSot/
l2KtemNRM6LXt7b7niFN7OhnE6/0dkPbTaC3a6hoTVH0ud3G57wG4cS5kmqUVa2k72k/LwMi3YZE
gbAqRenVR4v+p8Mr2HDLPlhA0ITB5edZoWt7oJE/21lzwXVyiCSwpigcCQ+ysJoJsAKa203rayvi
9/l2DT9bOevpp1KKG9LURTmODg5OAF3LfJ5cGY7PudB4L59a7qQ26mxPjEEugwYjecoWskyCKF8s
MTD8MWDuvF12o+gbT7I2nfqqRbP95XaUVOarmHd9P/rcM3XkApnmVN4PWSAdJNXXa9jNfjKqnY6L
2ijV1E5P1W7gQLR/thpvMSvCJInBG7iMaXSPhLAbFxfFIgvM4nPHjWDNtNT7zEkW+LIyzlZjshpb
LusQEbRA4jSqc9YF4Y8kUkPgSNJh1DJGT8NCwHvuiqXbJ8QTMa6A1W7f8Ff7nkh2LGyRgR3Tp9ar
15qtxL4vCloR0qcwyYpYEMPeDi1poJvsq1DTYfyeXPJCtAZcowss1KtMYpf2uk8pLPu+O75pQ2Ce
RH53imFZICvoqs2Ou//AsDz4yS8SXFK/9OMAtSyOT6pP5jqyanhlb4kevhy+5AzUoGxlOUvP60C2
podb5LsK1dkvJtScrFb1X81lQkPRmu1UCafOOk8FsV5+x9UeGTtSIfcI1Jrp9f4xOMY9cXvKTl59
exYCSN7tbeKnzMUuyLXjhV6GQFDb+Yho+Z9LyGKbr9prX4ZBdi8iQLrpPrJDd222SiwUNrr+W5WU
tcJhc4NmhZ58/n7fqQlmU9F1JxIzYf5mqCg4gedZjZUBeH0NM8MTzhXiK9MOkzOglZ2si89VL/YN
O06tWxowus1wfuaD9ZiLdvNosHhbkYPbir18QQj4yJonYYrCAy0kYtzae9lYndFkmbq4CcfUmSzM
sUijLedSDYYK4fLbq8Tqjlsu3WZCHeTcZakvUIE0H/d9osOOj5Eji7q34rr47jsngLE/C6SKdhYD
eomjx1q5xb9MALwhsdoxPQY+CF1Smo3GFrJvNoNSHY17QPK7o5QhSlb5O4OaR06Djv/fHunWYl8T
BBkCUeqexx3tV9LZh/pn++f80Cfv7x08Y72XiTLvUDRd+dmNU/Pu5fgp2TKrjOrcbzV1+Wp+kUUA
7QiRIwlGyes0ymgg/AId6H2tcy9WkpsGgbjKc0ZJZCiqzjmqWck4L2H4u2dRiwXZYqc+bnh6m/tl
vW7xQ5K03KgBvIk635ek6ImD9nqi2Mh9ZAWlczi72tVBy1EOtO/JVZFs+gBiIcnRz9WAR19+ju27
15hL55qvI7ftQ/2UrI++yNNuNtVJALFmDpLincCi4ovbSjHGhkPYVZ2seBUEPxFXl/yln3z47wTV
Y/oEarsG/kfThCsPwF1MYodI6IGwVtAvqFOQJRFkY5f1MMc/5TuGqz9nnLHiXuSo2QIlv4xHOGyf
+B5esDWlzGJ1bjDG8sahWpGCRPrpio3FLd4+iemooJePrl0OHquFoOlH54biXuiu9oQOrXoaFrai
VzGf80/szkuwZM+pwDiC/i7YStthcFCeNTzIdH+IzzLCbRcbDDRDCP48w0HA+wfz+D4utZuusGp5
CaSgfaHEOiMGmBax0Zk1u9hXxNT2HmST8FNIqz8gmWD3VqKA8PGEBQazJ4hH95AWmQGetDJh97zd
m6tQO+cntkJ/yc2qfz3jkdXg/K8NwD1+Jr5RxDFgdIcpkSNV8d88Xqc+jq2RBvj2bfTerYoZAjHD
ol4ADKaRszD2lOQE29kShYYJtpTFtqy9NZ/hbbuHO61+wFe3O23mgFxk0+zaWMR47rwuDqKdAd0z
G4IvgEy86WlIOyXf51eBd2tWhN9c3+Nxl7J9M6N/Idum3SS4cxxEd47aPtSLJ6ncaCPkUVHu20mu
Ov4AfhPVYVgUDT331x+gHUY0moTD3npzPigwRdoe7AAPiM3kOkvjNG4bmLIGI6iPdSXa0Ql++ZVn
/NeVZ9s0qoCNL1iqwRJpM8erBmv/1fZYglTJd5fG3eaM4kBki/yEFFF57d7VA9aR7VHf8WvuDIKJ
84xY0XVb9UZgwESTwI5zNk4D5niKR5T6cD1n/lfkidJ15YPEaTMrJ5P0yaQtlvhkNLj/GGHMSYFc
WTi3usna4q2Q95TXsZf+9S7aPTUBpzAZUqJ3XXGcQnsPjAhtvngcpZBGZQc9B+/pHyjqVJvQHbCZ
zE95fv2DO/2qciF8XV4lqfslagW/ZFTYyzsbwSPX+/SCBEhussxvM5XUCD3a3mceudd3NKWhG7Uy
45YM6DW/X66xtyVv9R3KR3OEtS7u/7m5PI1LOybq5MyBJDAdYGWF2rckXtesr1dh0Lc4WkUs0yop
klWQqJbPcJbdOfLKpA4aCfxBloBkfIzyg4iLlR7qdLotCbzZntAdT9bsktMcZHNAxmwCln+tVZI5
iwNa5UT3aLhplIuxwEdqVr8YxuqoMattBrMMtx86kg6ZMJG/s80qmMYK2UJSuszrBERfff/N5+HU
Pjc6KXdHSCsd9MVkzQ6dSyXAXOj+SD3eURlFQ/YSPKePgbH/ahvO3xxYJs8nbY71tZePoFYJHwss
RALUCAh31O5GGfuO11A//ZzKKZC1vKbeeS+p0mTjj91UzgSt48w7dq+urZE1JrYFkklOkbrB5mw+
qQJ2OaleqiPNEqrtg9UEg2VHOQIgBJemIQ5Q4pDC6LRcz7nUBjDBqokR5iGIecikFc4jf72OF8/Q
azzYuC3n0T0vGkeylZ6w7dRdplYtsgMtcmKXFqhWB+meRRzeyH897A9wTkkfsutejUvETF18Ik+y
2CirZyPpj9us0MD9TtnDroXO4/UIx9sqhhkak2eAsvj7OiurOCOAsKi+ml34dVBeGZVivVTad4vC
f5daGYDZd3zGEdejWVEbbQhPg6lalng2RUGo8cvbhdcxJHknMG69yO1CXtOLXlbdi9ojvkeDXR7o
6yfuIx3n1gUh74ToEyyZejZAj9Bw+3aqICDyfO4j7tYcTzc1G6EuYOBc8F6NOoRhn1AGkuGiwt/S
2W/OhHxQzI8D7uKCIVnmCjHFAyf8Blv6g5VaGAy8KSAVWAG5B+NOtp5ygTPE262P/kH8x2Cj+1xP
tAecBSrd28+T97W16QrNzN3SB4xLwVol3q6845gtGDPJI0NeglBAyuNMnIb9nXccgQaJEUPUV4xf
fOxvBSfygEUmi6aFZEo+eFsVC47TjZdYH17JgDQlK8oQ56L6O4xj/0XRW1qfMcb1GjVXAtESMnmR
tGQBBuUUUiGz9LfJCdvslAs1C67olwMIboz3zE8/YEIZvdSQcMq6LqwZ9Gy8s/MRrgD4S7IgeZSj
51Jy7+hzotPdyRnYlFqs5tQ4RPuIG94Ix3K10N0RNSW5xrcTPamqQvNk5DEFiY4DntXAUQExMgJ5
PpOMfsU/NtaoNs6V5maVgo1vYOO4r0TfvONKtLxHpJIFJiXUhPaLtwyky501NYjWgKchBwpPTZ6D
shfk3Zwr4QVMLojSZiharGMW0aYRqPzJmYTPteVgU4sf6x8ufrs+E0ECKa2BvqZZAahdTElt9me8
LnfF90dLIsbBImrUYS8dSp0UCeVJZ7bCccGpy5TsvSNUKw9V51llCS5kk/m/FNVzdvUhJe0OsINv
QP4qgco2LZrjYl627eKXbSE1rdk5+5Dg+S9xQcIXWnWu31DN4f2s8Xq6sM7vIiRBgS4KitE9JRSr
B1YUgLY8qVUo0Bur1sQO0VcdtyEIt+X34Z13fJvWIXoNwM1/fZmPDPxtX/aoYI7WIiFvCDP5DmbX
qrYLMkEC+4R3ESERfzQjwEqn48dNr1ihS90NexrofiRJ2AuYcCA11pO2vyPWR8f57FOvVB8v985+
egU3+QqDxYWJWQNU5PTxtw2j539N1Hy+djmBGEwcr7Fd5LbRedvb6lPI+QlImHp5FIYMTl2KuJI8
tufLikkczQXliUWpBfaVMg3nXVRmclr+t4leNos2tZPbvl5GpVEA2D7wFUpzfCy+iNWl3uxc66qY
6kEPQomVGLQebAhgaLWEx3g8QrjYRoB73A8hPkZy3HITggIQ0b8LUhChjx5SL5a+OCt8cQuZ4uf2
LdfWGEB1NRJWaW05AZpz6aBYAX1Tdv1MYOAnRNomtPnJcn3jQMoooB8CTh9ux8mCwjrjhRb94lIq
fGokawcvD5GTuaBTVl3f7E3Ln/TSXkcN0gUVUfcNsMG6BeiPimLKnUyk8WESKhzIJ51pZYUAMZ1T
Zf2vsR0RGqBF50Yzym0jV4cg5ekUXpoTB4myi92d3+wVO212u8K6TPiF+lykna2CTAmOhNGHwwSS
yA/z/0QhXctF9jFkAIsdZ8Gp6XebJPuTtPhg+o89D8G1e0eFshFeHXkq2vC4/1oDOHTSoXQYptro
hn+oEczH3Y0CP6akmT41b4XMMSpRiseT4BBvm5q4XJjEyYHngUzHWd2gcGVwGX23Ej9fGmOe3Fs6
FftI+ssrcrxSAGuBbtugp2EdquDDvU+2GYBRQUw5D94QhIueoRXfjauC2tIBeDfJJMqtSwLRNF4F
wWi0xicLFa36UtK9aSgitOlyqbCQk7encbYDwZ6tnxWI0AoYM/KTy3OlW0Eib7hjo9cj6nbhsrPB
q+bLa1qU3+wGEeIpl/lSOCyS+svg6PgaNNKLapjD2kjO+8cpUKpL6DWiPhLvA022CiXTrr+aJQ5h
Lq7PS6szwAQ4JoRHfGOy91BpniL/ZMhv5i0VU98xGAZi9JpJN/c+RhCzocZSuAUwrnZIdYaNv6+M
pcfFCs9wZVKjsYtfH0stYvXZwTqYseJ4NJt26gubgVRFF8u07XT40JGKqaiEbz7p3vwMGvMJx6D3
bsxVj3qPcK8pQKxCpYYC8BWgF+pvvN/cBCuJkz4NVrD1TszXGPTU+2N69rZuu6hXp9XV9D9/PJjV
lN9mKZW8CR4CdhMGVYCBhIzkw4hc0L/Ejtx4d1EkOrkcp5+bCSUoaQOrv9hvnKoqS1vzwNSumqAN
uSGdRVJoOzMnQVg5l5moRyIbknbaUFKL6UmuCexa94npMrrEvIEc6w7bttx95RaC3nm7cbe+uAGC
acpT2wVGxBAscpvydcZh6T2Wetr1MQh50PHqwOxAs9UGbYMcd6XAo2F+sKrem8PZsgITCvtEguEH
RKD/+UoexpJqMatcotzg8kRxCU0VrBSrSznHNvRn4YrvbTWCPMan89CJ3KZH0Xtkt2QnpxJOm5Xh
vYuZUvx1sxEmSZ3yP1bTIRAqa9C9lbo4E0hZjmy3ID4FleQq1aWjxXXG5nOTDm2TtpzibYZONaeG
1RBDCONIPVOQ3PII3YFK0089ASU/veQfDVEntlNoRooPHRMbLWf7JDv4RSl2iqflRvz5HrRFTG0R
4uf0Ob3EYlM7U1pTVFyx2YYDLc7hK9xej7sR4pE6qt7u7MPFJlgikYv+DQOCrHYqp2DEa3Us83KM
M+Rzls7iGnktPFOgWEsasnYvlsi/rRtXaZBYA+2jXrYvV1uYSmdPokYh9EJyCXSqtD1r+ZyRexTu
MXilEKhjcfkneXSAeA8XbvxhJBqyIJZHXGkJ72ACdS4Re9nL3X14t/82cYAliipFcyvrWz/gX1tQ
K3xYvdWRCCdSAjqxBm2EFgQl01Gi7/9bKYXDWasqM381OWIhal6lhzg1sIaTilT4R3LbCSG1uuFi
wKa9unQqEueOqjMFV8YDgz7Aw+PpMlXsl2V/QTedWvyi1UdmfM8UuXr032rtyGi36BuUL8Jyu+Yr
nBSOLTg+yfOW+ytAS+mAxk/rzp9Cpzw+b2waHXo5n+EuNUeRvj+qBDL7u4EKstC1N74b41qI05Lt
TX31/yBQUdcCLdj0y7WIp4+wiH2leBMM846SadA2/suq7SjbVE/OhH9A3GGU1hXPBMElFAS1LLsk
mYvacoSvjw9b3eaYH3KzJjKAFefjHnAc5IzkSvypyKZZkTUz9VSOKA4gGDXXEBqRpYH/h5iZc45A
yRxlURzQN2HG12ebfsjNcnhEpzeSs4QuuxC+Kh8WrKrGS8XdNou87kCSWtf9wvll+8SVct831HVo
HJJeXCl714if3Kzeso0cZphaZvjgiAfcL4AzMKe8NA/XdSX1NKf4Tt/n28bdBtLvE2VpvkWlW7uh
Rhs7/7d81EMd3vrZf3VEi4WHBC8/SyKxqCJ6HOsc2ghr52n2nXXzWwJOfbvHxFP7k5xTM9vVM0zD
AROUqMxumK6tdIrkwzettrwhZBJccXbxi7LHdXCHx8Q3G+4oLKr5Ou78GmDUy/rxATJksc/TitC6
tTOXWYdxLq1O03j1HfkNelqKeMHwLetILZorED6jpXYCHqrv4BQjAmbtCsDF9dH3bayb3no0bHQE
qbJuBNPATBu6pt7MPZ8/yNeXXDB0qQaRoZ6nX+X7YUK9PpHU713RzfMoBljrZpwAqKBUYxRG5MXJ
OHRMQnV3KTcpa93iQ73a0E7swgXf+R6BiH/6QKyyv8bgsmzT/UDIMT9PcpSGaCtA37XXQ63fajLs
G42ORAnFmuanQDxkn5UwY36XDQ2E5kbzHyjB5dc70/WCBdKCrR3LQsebc1OXTVr2RhSGAr7c+4rW
epenL8ryEPRUg4JT48enzBznMWmy2/xbnqrUNu7uE81eLt8OeelXj4qH9jhrRx+B3u+mquOFSunK
qGGwcKIZ7ZaXtsN/wFRp5gSmoqGRzDpp/LOXzYaG5NklX5UeFWapk2LTRqz4SwqIfBv5UxrkIG23
uqDCjw2K93vbzeP6SpKzuiZWtxYYCkH5vB0Fe4MOIYVX2/4ZGPHEj3FVoWDtNiC8YbtrDxXDCKq3
ans6ariPS3EFN8YUL7ENpWYY30RKh0o52AzhrZdPT6yLgG4rGqQnie1zEKTaeFzumk4nedBwzz/h
h0eGYnGatLjspaKwOQbsJlReY5af1V86xucdI9uEwUj10c2ipP+jef6o7Yo0lrBGJhBhJ/pVPN19
aexPWmvg6hoR3rBgcZVWSs4bOqI4lZE6oMzanPq1s+X+NJbXOXQ25pSTpWT7FolGK6A6JwIh+AT+
3/cDCnv+1gOtNCnSboxdAHkkwQTlQ5z7OYKKLRVS0twaKvuPTmcJ1I3WSYXCdhVVGpRXLr/jZZRk
pTNhsBQpxWgEB3U8YAX2A6m5Z4s9U8DhXzsPf7Zvl2M0C0Ipg1evjjAKOplB3IR5/+LQ+YlBxkwc
YZ27WwaD40oauUx9LqRL2/aXK303pemfdpiMtSLCxiZkNf8ZC9JSdlUP2OQXW5w+bS2zFssGm97d
hPk3crst4MxJ1ywuqSkV33VF9L0ku+UW755GsBNXutg/90icWGrB6PZrAmSNlNtwJPC1cCZa9HhB
vuVIAJ66zrE1nP+Mu7h3FJkyhOJDtvvcnYHTG5GXq5tS7SIc5DG7dD5aVRKfGUoqtJv5AhxyO2ot
BQ0TcO5Vi4FxepXmRoKuYD15yMhzyZjms1QkDDRStgDdZhSh3Y8NOLQcqZJ7ip+Fg5pI3lMM3sKJ
aEftB+JGvSpBhKMNI1Ochmrk/kIiUnjkVtqEJAHfnE6ZGHJPi06sdZx7H2rhmAyn0pFwIF3pkCQC
m5Qs0Pf0JxvbVFZFrEMxarfT92BCGVlKmbLi806ONE8tpVDOAH/GuP1kDul1d3xPX6JdsCqf1Mfl
5kminn9dA6Rw/fR9ax8qvwUGH9miSXrFUTrjS1VI3Qu3Y3Klro3b6koWCadxOibcqJ+/1RSGO1W1
EBig3E5pJW3ve7DukIlHZw5/WM+lLvFexpf7/oODSgdrbENfB49H0vPd6Fe08mPUkRAGgyMmTHPX
q3Y81hdFduMDiLNm/Ka4yO4bl6ajQ8c8Lspv1ekI4JZzMUyxva86t4cxIuPXEj81IpFldycMe+1p
P3zAg7e/i6TdIMWH9IEzrrQ8yZiGKgKTM9jrNFVnkyR9ROqX3o79LPubcdzLM8QqZTa1niBOG8CV
nB4EbSH10doBufAtqtUiCtABOcNeQRNonTerP08OxHgQTY3BsFkoN9dVRoIrK1xlyHCxL2++VEaB
IVrj10MSROigwFQ48Ve/bwxy0BqeBwTgM6f1kxMgAfgeh4o9j6t6TOfX2xH+MPTGP3DhH5LkcWbu
RxTB2dmc0EZ+gOTbwYnKbSs4xrUnGG00x+ojdGcUhy46KPxaxUv5gAD7juKii4PbXS3kiO6sS6KQ
BQ0yrA0/lGYdtv7H5eDft4AAP4fE/Lz0f8ZaTEcbaPgKsbcd/TLajnueubKTxsWxAdDTB+jszTR1
LvzLBGuzftZOb+XH10mAP3qISTwb80x8NtndBzl7IKVAm8S0udqcMRjSi4jSs43F7Ka11+dvbsdp
/GHNAjWbROUHfCvpcNDWyKQPd8R/UrDV2TnuSXSTmwb+2Tcmaw+v6QGQ8fBx25Pa6PUI/y8z7oJ7
Hptlum34bFX7Z9NKpTd6+lS+pSbjRMlNTQy+ecaB4+r1RVVl7dyA5xpXBIhIQFgccnnMxk6sPt2C
y6hQhpf/iLqtFb5eaNMgcf03P16owSyUzVan+btE0AdTrm8bRcw0OVBSzFAWWTY3jQN7JqvSoq4P
altsBzc3nrscj0M0XBNyArB9M5NEnbcUJKBGt6PFzAaxSw6uQnFRv0JhK1Oo4fgGagd/9csHU5ki
vXk9rABKmc8pc7ZJW8O5Ynra0tYzMI9vUV3QkMqwjY2H/cr+hU6NyVEgZ6LVnNMwnTBw8QK1mZRk
Als+rL2PYr7hyoqhFRqKmNGeNO0iF1Rs7RSewA+S9gKqm216gudjL/pCgEC1YkYX845lP8YVgGsd
g4tdhlvy0xHrmTQvTo+lY81AzCAwkKJJ5CfZ1pTWm0hf44+4ktXTg+hmhouDWvHkP1Gc4rmZlDd2
34vHX31gWiTHZDAga3maIG7ixtSSIn0Q8HJJT3/awIxygdVtf0YpahUlOQzJAJC3DzNXUpq/raa2
0XbxHHvMt3KRL7iFQtveL691cjf5RanJBHonDhebkqHS5s8bTqpU6hedwkF8PnZlev8amYFz6yYl
rLxrkRep+gpjMzwhC6/CRtrpGrk1LI7pPLSU1t6wSyQwTB3UdEYq1gcSQUfcmosXRWnw7OkxPvbL
WPwx/qxPnrONgl0qDp7GgcMc3YzTpSK/At5ZunixKD6T3+SRrXKyUxJUzVAO2Act594AF7vgzsP/
D6sfa4UK/ucAPKSOyr9XmN4AcAH48/jyQix/XP6Vo+H97ii2nyELah0Zeo5eKduS8nSQmK1MphIP
FUHzEHutN5gQp0zTUog9j2Pf2QldWmETIUSi+0WKQF2GPOVE89TbRktE+LyYqgfp3uqHgog/UBJJ
Vpv8v9gHEDCufqirNXODJ2hH18rJVWUkS2uKc8pgKHoUuIdVMoEXWq0jkiSIMLKvW1S6WrQBRH+z
f9PhHiNA1AkuGHkzLMqbN4511GlNPXZy4CzS2oSJSWAu/of7F/MlplXxLte28FRfdUEyO172yEZ4
YrtW3JvvX6dMCPg7fwupzYG0mCKAnq4Ad+xoDMjClqD55F08Uzr4m6WcfAlN/DVwD79Y0paFIFvA
qSulKuS+IlQgu24+DlyJzD0zqcYdQvMI4v99m2fxHAu2yHjaOs1RYSOlTLB/Z+eBKMe/ZjVH7TfO
/W8M4ouPR8aSZxjpkqZRpGDgSDLRObzshVJGQ4G0aOUyfYx3JmLr2G/5k4/DfURlOaoedysFV6Sy
3aMAZ+cILoZTJz65OFaP7r5bH6netzMG5VolZrh07nHlzpwD62bG60co37q+Ajd+bWt/uquoaBbL
sE1iZAMR4NCH0GKPFE9N/77iwK7FV4IS5sMwnbCbzpLyx3EBCR3xgIF22HIZMzT+j9Jw982oMIWd
M0K/fSPdzJXd7KyGMtJqGKelpEmOwXDAP6sjyoTSONy8rRWP+IJ0PlNWK58BODDNOMwEchgGY17s
L4pqy8UJ8gNqL1XR4fjspMi4x3ISYspSgUXBcRJnzXzHDV57RKSKBa49PamU6PEe+J61NyuA53+6
d57wB2nuy26Lmj0gP6c+9h7tY4GL4rc1O+/7JuiToW8VGRXtPvII7DtsG1Womao3ZmPVC2WFWtpj
LZgzBJXVSZOo/lksAKlUZtcmTGrMO79P8xXtYi8nIogpz/+CFabicZ90X94WxdJPLt+EnRAxYHjA
NTj2hJQJJcJS3115BhhpEIYqxCxJKyZ3hvtLK16n0/bgFW/jrM8n6MhJ5O6BrPSF7U7VfO1zR9V7
8Z38trRSMhF+mAODF28gVmOAZOJCDhN1aYDiYl9k5scnKy75EhixfTErM9lnk3nVJ+X4059ui6iF
z4heDlg+8lTtfKkty96325qo1HxGxxnoLlQPZ9T0bHuDpIUPYQ3WurPZhJxZXCovjDCCB3PKm62P
A4YK+MViLLPROllJoJbbnEHK5tS9S69+uvTmZXuy/kmY8X6kOy2KSt7CbqaCJ3J7IrK8oijWKWsh
bazxR7po5NkRC/wSb8WNfUsDmCQrcACTMaxdHeLUEB9fIuu86EwBc21oH0618IFGj2yYU80aDYua
IWGKWBL4va6DEtlsIl4TqmYndULnk1EITIXtl+c87nPtA3I/fse2fvd8hISRU/Js+orFCn5UFfW2
GH1Z/Pom2YEpYL77WJGKs1LlMZBNhONOqmqPVraYxClje+z6d/FqGDj+V7uyFdFILeGILvua925F
jW04WaeBmewvhNuoQnQbx+ZJKqllJWGockI3g1sRr+5fAlsBey70sGi4+TeGz+RsnKkaM7hEfNOg
DlFysHtS9FNl7MKCUqsJk/s6VK8YoN7sTe+iGOvBeL0xhgIYFZOXJBMyMxPD50oODBjb0ylkJJYl
RgHP5T9ruqTfEi3fRkSXWoNOjAETOeeRyarUIPnOfzaeli7HR2cd4eQeAVuMPMxwk1nny9+8KS2I
kLxVkOinlaVvQ9JVT2zWuOjM8botMgPD8IlXIQRVrorD65dYlrLClLNAJt651PwzkANcK6w2+BbZ
QcCfEkbm8cK/MiytpwJLjZv7WvrAeB99b5igHC0UVd8xRnuL2FyjWM32VF1AdmrD7JHN1KXmrtQo
wcBzd2BQPb3DdzSoVoLI73DyW4+RmcLw3qrW7wrMYn37+qF71bxS3Qk6JM8bVz+64r3Y1trjEyZb
dXCxiAYRYaQL8+A7kiMa0ae9rNKyyuRi7qU57fYBF8vR9nZUWseGfHlMe4tuX3HJTS3+c4Dcz0rz
oCH/G0PvrgAaYENNmt1MFHpnq6Qgv1gV0z0SH+KNNeT1L51B8Q9KZnkqq8uWotgpnA7x2sLf5400
JSrwUb1V0w6mIvhycElyVltqmv3RKWWG+oaaugaLt9uJqnArFbenJKmfPZwEeZxQcWj+1MebWNZA
HOtHb/eyp9LKX2H3xYwpbO54iXKJjmD5bjBlfwa0L2leylv8+smwDDEX7/9vK4aM5ApLTxa2t6/t
HYNEDPPcin4N/wkiWHQtwsRNu19vmImsoM6X0pdtywNVt7EQ+WjPSNDazKyGh1XZJ1dOiHz/5p/e
Pc8TaZ8SjLZvSKo/yszBOzlYiUKA6yYHzryDyX47SErpm2ZAP3UzwwJeQcafG/CGj37Q+yCEJDZ6
wyR8LjhrW7o0YkIlpdbXDFy9r8nFvOy6bhaiPD6PDlxHbtSL5hm/GLrM9teYfduTTl0XRR63qKr7
C5vPU1hbH9BxdggOiEmDYtqQM2/kXzN7Dy5yHp5EY2Bz0lUPWc27husXBYx3x4K6XKfza+GdKdGf
vHGjtwOSCeQO3qWPJm7Pruxeyce2biA2dVMPCmoH/aC6Hsz+CBEjoT0uvQ6R2bYK0A9gOv2k/5mv
yIrc2okUf+v5uUetE+yVTfpza0ONpNZRh6JWNI/7NHKit1r+XIXgHE814qbfrSfz1331OOWBbTz+
5jdrLst4aGgLOlirhIwcZ+qwsALJ0VfI+76FVTv67fyn1yD1i9R395oYcpkfGcto2bj8HjadG8bN
u18SyDAcKujgjTm023hrjUCVll1C+6cCVODdpb9/ILXAel7Qg1SSq4disyn7/jx257D7/LtGyzOY
WPnB6C4pR4O9GZ0oxPh3XNHQlo6hZ4dmUtSgqd/PJ52g7/Psy+EUs7YwzGG8iElPtjLIoueYBEX5
/Wq9QD2kPYJiLSR3ItiWp7edZ2V26NQkvzPkN1wtppRckBRMCW41x0SBAV4Zaa9aVIyJ7FV+n3zW
Jj9a+YKyOpOFoQ0+i8xsSyw9i7DJ7DJ9MF0UZWCvPxS5LbQ66u2+jjCMq8+Bp2DvywU/Z+7sM83d
Ul+joX6s5qR9oMBD/EIOaujn+RXIayVgZQirig+qXNAh0zISSWct26sGCcS4R4Jq1+FIVJiI9lgk
9r/u7vojD1/R2cG2GT8Zeb4S9OJJ0rlOSQULW0tg5l9ybeJ+1AIT2gFQBBezEiMUfAhfx0HfWiNM
Z3fzZjpWYgDv6TldqLDwcTAZpaVY0y/z2DZuN5F8nw0simh9YuTIb8VmcswKTFCD4Sc2rlw8Srws
P6j3a/byoFkbstEHrlDfDs6pkTdJZNZvscfIzNRjdKfn181z1KxaMKuVSnN9dqTAEANWs7VDgjbf
pWYQE9nKd41rBLUWlcymqXPmjha36u1mXlKdhQy9QsxVJAwLCcq23x1hS77Xbo7zgUd6rkz//7Zh
+5Mr12on1EWsSZcNDZhYpDM5fLswZsjqAdPGiQUewhOsZHsSA6C66KgYVXpGZ3vXdIGyjiyX7Im0
I87yVfbTi05AQlV85Bf194IlStjgU62ikEwKP5MfY1ovg6jZajU0/5n9SN2r9Pu26/VfKtsThsiG
8JLXCCEomHvF2UlMqLJ6CC31nExoA8qOnw6LUmhINQP4/JR6kszumUs5rYDAlb5RHjaQwU5x1VXU
WPCih19Jv5Ygu+UFmTw4pZ/DGUvZxpjiMdHWMFK+sh2b81WVhwephXV27Ub8Lk8/Apd5SwYtpTtl
PNJHOO4ec84WuodSjbgHmafcObSK0cqCldQapBXpC1xwf934/Nr+oxtXVn9Dmp8pfsyal0hZQX1V
S5WLhjjH4gDmrc4i8I3VZ3bamD5pI4P7lkpSvJ7/0PoedLZxH1yEs+SoKANn9lq4A4l56vjIQTmt
S5J4JdqogNivYxOzJAgOfBrPjj20ZM1No7rQ6z2ejQS/4PDj+Z3cspK6PsZD2Qn7mfGM7FP+4E5G
MDPNB3ygdWCa1wjIudLOchIKNNQ+2SYmJ+pTz+2ClQxAnNQjo3I41zE788nerQ0fuJWiMpao+e/B
7EIAGQB2yU/3nVHIzwrMP7RAToovgxN8CAmTIVisNukyhiTBHo4YZu/32eC3Ar5YK+UQ9gtjpVgZ
pkqkM27lDzmZ0hKx0xc02zjCoeG4LamPsNgz6K52EaJcYySZ1uL3s8MFJIsvMs0EJI3JsotesevZ
cSTMz3bclACntZixld6ZBktfuGMG2UGQgSW53ix3ORtKJvf7JPZr7HZNqTc5oB30LVqqZB/S5Ykk
SjZYL4w5J//Rj7B8Z7pgcER1HQWaAG4NHF0WdRkz2B7f37vrwc+Vu+MMSTkC8yzp60o99r0UQogs
NiLbosNatkZZ+mjvrXlLB5zvNK+Vz/HcjcvtRN4P5YaMhYN+V91UGppmh7KDyo8usxk1A6v8MhT+
hP2vQ6c0aROplaNXrOLM3re5w8gOyZO1hMWL8i/grZU5W05zokYFH/QNY6MbtXe1ZRuLa/V7p8rY
I4dDxJf5okw44uqzvtvRfvFQuUX0wbX1t/1MrDR69ybhk/CMv1ta7CgypzgKKrMmCUb7Qf8xt9ad
BBgLAKrU3ooLLPwyAivUZxwkxWBASSRFS+/pQHquMXj16xHkZBdbZPnezzAWYqKjR79ncc3uTA2t
Pf1KCWENCQsOVr78wkDfS46NuMT4u75u4ba/ZTTbfuxwHSpYlghUh8TMktExeDJPpTsFs7W279ef
tF55cEADpbQLoBZN4zNOo5uKWrXgc/8pW+mriXpwYUe7fIY1F66eLi0ofaZaBREocBtachGpApSQ
Mux+84UNSPC3V62W35Gk0U7/FlY3MirXiL35s8rRC3qJxKkKS3xlipWj48eFQrVdkZ+XIcI6RFNu
qu9t5jJLT3WjhPoQwCaEG8FdJZR6J33LO4011lFH13yyQDxoGJZjpvH99viuM//cCBll4IuaZvXb
ajBrelWBu63E2qSKEZS7zAl2N9p0UibwmpxVHC4Kfry+lWZuShNZfCSRp7U5/srr0OAxeic9e/ZQ
QlHL7CAq5pu4BtDskmb/NXYVY9TAGya2DgaTU7lUUFRwg7EVh76TDPZSMKbTDAkaq8dxosFYcsTJ
4q9h/yQ7QnOhXDqUtRhWsnDVwxZ+z3a/hWAmtcPSb+JyrF+AFi76zl+//eL8rrBItuhn369OICz8
sYloIKxdTSvG+Y4PeYZhjiidnxNPsHl9u2P1Fl2txdb9oMuZoXD53JPF9CdwClxDcgcI2wdbtO9I
LLzL5AVW39GfrbFWdPGkctOlFTCfqt2RznrixWvNTsa1VP4DfkuREdMJF2ijuzJ4Un0vQozW4EZn
5N+MZxv7NxPlEyEjJwPPh1cRQZ0afggfAUz74YFcHIE3vLA1ouOtfqwqNLjdd8RrZbMbPt1J6ww3
x1DF7Y219K00c28rnJYr2iPpPJJ+4eOgcQJAgU/uAAw+zFUl4SVwdPrri4BBJqdpNydOLugWTNlf
doL2mO2ViV6EyTwaKmBt6MPLq3hOJTRcbq0zrrM0UsjzNFFz3eAQCOLo2FahKn79AP/G88R2HWLm
gyuitYIIuscYhKTALDrsFzOX6wttgEfgCEkDTJolUvqyIxgIiPzpI0u9T3PFzb/vh+27KLN1q1PV
w3ECQwLJxNXwMAlawOo0rOCIXlbfpV4VD0nFmF2dTKxT1DPT+Jn76lJxNoVqql7XC0A1YBQbPbPu
tNrp3EdnKWQDqmwnlr04gH6fXBxuWfV6LKbwngIDj8fBh3yjN5RyD775KpQGWqFN1wb/euVvKaRO
6z04od46Pntnyof1A75SwXuR5fpHIpHshRT1Yz5B1mCUjgc8pcfAiONQs67hVilg4nzBxgQSTGpG
ydwesHJg8UpBfic2b9ZCxNMiuqsWmOB3CnTXDyynvUVBfLP/JaAivYIDDErQ8KSBx1dEQyxzn421
pdFV+snLc1HEg/TpdUlJlCyZV0JFML8qocm5h+okhkkaTKti3LXLalVdy1YXRxOvRgunaZ+2J0og
4dLfbNxFM3NGme1ew9qYFNCNhWguPPAHwE4OcjDM3AzoBTrgimykNeh3ioglYImajP5bq+zDd/Az
iY7SWC/czwCwRPar7uCXwO04DP8mAozfLWeHAYkzkcsV394c/Np+L6hp4Hpet56MsRB325ldom5e
72no6xDAH3BdllegizOUlshNAll8k+xeLIvnbFgua/jpIQBcJU+Bcw536adUeKokRtqCvNaAri8h
EglKNOKev7CFXweejEJKvqu/3s+S4Sdy6Fjn3HV8V8H70q7Asq9oQ57g8pS8ZtH7bcOoJw7or8Jl
cToPJxhPUfa5U+cu379GUkWylm38qi51HwFK4V1boY+oSLOjYoX9kpi2/73TGmaroDdDKDAI4Lfa
fFNNm8kyX9fgrSFNxBzfRAxxO5KlZ7XCOv6Ks3lP+PtWzQmtKf7L47rKp1ljuJlqc8AWVJU9EFAm
TdVxNBHdhJL04Md74GjMoY1ViFa8GkXC8UaxKjv7mi69lvZG2CmAtZhjjxgSXg8Yj45rdrdIxAug
B5qR6FzHJSs76qOyL+oQQwQF2Vp+OThIo09r8WOEGlhKdxxqtoRmi3/gVXQV6qrRaxEuvKHfn4FV
Jw8kmuu2Uq9JhYpsr4xrQPG6cQQSdGDO23CX3rQyDX6WM3pRhzfbgVDPT79ioEDdivg9nTAIMiBk
nmFo3HTSytviL71BkdkHCmm9mV4ikpt6unw3qaMHdpNeeofwWhDEbKKUpBdAd3t6c4A4rubNyo8e
jSHqBAtPOl+jLmd5r9GqhwtWuozQNn9+GUNKbkvIJYL/GMckBKEyN5NiquyRAmavnlDjISDMBCEN
TPdAjrjyNm8q1Qu1RxhVc58KK0UXfSEnMaKZ2uTD4A99D0V4KKj6ptlbdH11GMi5Rir2FuW0I2Sp
DinAC3mRQ1VDvyvu9N3MClGkBN2W1fOU3ecVE3ZljclDV7RUzQfs6or54bDXjVyaTKa4PnRk3sRp
cNJsYoogR00QnmAVwWEKDjJvmP3uVbZ9DLK66J1XrmMzZ8PhtVzgmJLCJJtVvBetbDy2sXyoTyCs
lHslwJGY1RmyW3M26qTbEh4qX9aaQFprdVkVPc7DT/Yp0U0iLMT8u0xVPBlaeY+Gxa9zU2jLUNiw
fOrS9CVifZhOweB2PhvtKB0hUYboZqEGxPnhbTR8ZIEYLnPuv5Q2TllHgaLEXfLiiAK1b7/O9mRk
t7jyfDqSuaGU+hw3bH8p1YU+EDtBDIRv+M4FGGR1p27DX92H3cyi+Dj1CF6Tny3qa2XDkloziph3
M3c9voloIOV6Cejxjc4X+d+80ZEliObk0m5w7g36OUW/v35+TiDusvduuloCWZsXOoQJaD9qjR2M
sDHxQx0+PZcz9HeL3/7HYbWOI1IL1qXMTUumzFTZIlmx7vw31Kj1IN56MNEv3N2PDWW8fiLpuLFJ
s8KGnZ7xpcrPh648dGsYmV90TVTAKw1mvqTIkICjm6DomDesRB9/CBP9OKSO3dREJWmb80p3UNXg
eP7u44UOlzLwcjSi+sJNrDHVJiO4xcH09bqePbL/kBqFkxf1YbGN0D9enArU6fTVeYZ+50DSdGxH
IXpW8TJMcit9yROfLx26B4Erdw/iwtFYUFtbW3SdpXgjt3sDc/Ew3gcvKBw5iepBcHb8zjUsd6hA
ugFf2pYw3OwAXJXVsxmC0jwtEFmsigrVnbgt6ogqTIYdzb28UpBTKYr8WE2cfJ2Jl7bpx6edos0h
jmWN3DasdetnAkUsZ2JUjNxxHCPyWl8I+hesGE7b7lN24GPYNQlaL3Nsq9i5L8rZmfAOXBYipcFm
5Epbp8VlLpjonLYh7zopADpCbCGJTYC9yWXq2Iv00zQMID8mArieENHRVeEzp9+BNwwplZlIXOs2
bJyiqG6agonUkd4exw+3c4EvQ7mS/Ss8yCETzIwSa0YIYd2Qr/Y1FloYYSuxhHO/q1uxYe6ddSOl
lKikCj7H46ZdqzEjFJSPHIIz5b2lP76nf8WtMtf/0/L5KWQ08gJyrCaY+A4m+YFtvZrPDgEYtH+S
97hcPNjhF/jESnSExqS0AVMDx/iNRCQAsNELUKuGFMu6vS8192eMMaamx9vVBCu6hvodFEX4Jwon
mFdiu3UK530saqTCK24j2SCTipLFw3c4Om+B79qkVh0AJc1SWzNnFLImXx8PySuaWWXiT03P6+ky
kQSnI8YNXXqKpuNTKoqtJxlawptZf9wIn1qWK4DDbFXn7OAmj5/jCmchUnBSVoFql/QMSge1obiH
niEgNtqcNn7sNSTsUDZCGHZPogyfPXF7XOvf/QhpWGCrGEtVHQt0rJPxBjmGc9FkTmxOTPAFJ+Br
P+YQyIOk2TdQQV2zB0DyQXzSV0ssRo/a9qFRS2kdluco6ej6acanTAtvSg0+EEqu0QFQtOTHtg7m
2Lzw82ab01DhDTrVt+vlLFIKvyBBbCM3PSCYCng6/9IafX+64k5r6q8xlf/kabzVqx5jftdHndNU
sRsq36ja+HDDkmUO7uXv1D7DmADepiKd7lfo+nbFFyNsVZ2WjzOgF8ZZQA8KyjnMPFrpHOt9YQz1
Cj4ZxgFiPusP7ybEt4VKk05XxiyjDVrKircMs6IQBdLohJFY+iTeVfyhtmCXw52fYIzFq+paunap
izmkbyez9onzDZT2aJk2LRRMrIbMEIoALCdYWAJGR90vyALqp/XR95wDAk3MoZb8JDULAC9CT0Y1
N6rwGom4MSU9gnEGq5Hypsh2dFdFWQcAbiOaQ6D224OaphRCxS7EXdXUCgMUgVDM1kubZXa78cm4
8W+bpMlcblcwkJU7pTIsSGs7gcMALmFXcM1aD98OL2RRNNoPvW5dYm7quZHHsuJwx6Gine/aaHQ/
1MTuzboesBcswIZBF47IFOt2RgQxJly5Dv4AxLkJn9t3hFWG0gN4+7hxpQ0DIpumklbkfPkT+2FW
PoX7ObwfmWHfmaVhqAkTd68YtGM+VLvcJ9aMh8ygxGouLBv/CL2JvdFmHpotEVWR26DFLHKO+JdW
Bp/2+D91lSDn00uL8J5UFg2c7wrtxH88+UW3wUSdCuUeEEWFAV8l3wcvDl61wEJ8Ogi8ZXD6PcP8
DOFsE0v49iuHlbcTlse81QyXDXflw5iYbCEWdppADmUA2Y0jv81HN9a28Yb6jhNDjLq/2F/Rx01T
WkASRi9n1xd+FNiPaiKdSlA1w5W26eK6yf5rfSo+Ext53OfGZzAEEed/Q5ucLfwn7hLsO5ObS3KM
RL6UZvFckXJp8WtUJOGQmP1WrwOd0iKjUzqNQajOEwgGsHzjOKtgBvrDtV0Zesg0N7yZq7+Msczl
1+zHguJ+tQtyWjH9wCRI/P6kReKCCei7D0AwVZWI2ctZcfXj/EJE1dFqZhw0UFeLMY2J0niFv9RM
WQAU0eNF+Hh54ShzlSsI7MyN5UzMewVCO1vckgH8b+af0hO3VvtRp+oDPZc42qiaKHDf9G1JVUAI
CcDHrXs7fGI6Cyx6k/bSbGSHAxgPZHM4NJtePp5ECDG+UUrlGID87knGHIse/JOESBbbszQxUtZz
ypI5Tt9dQsz5SIT4YXNVbDArC1YqBDzpMaAhJu6Pm8pQ4HxuCw19mZcCIGlzeuYNaZ6mKx7ULnr+
kbmneFwLQxL8aiS66EUy7RZ5EhDz+5uCHRNLLRiI1gblxtW90/QZtjtHSAwYuUVqBFdGTudNYLCi
CHieXQDERCDbY+vlGRsev9fZFnh6ENxIH8fywe1gn7vdlwuSzg/bN5yTf9AWRtXJNFssukANqTQe
u3GEc88EaB1jPAdNDPbBNJb0ai3ENGhFpw1sEAmVV5nHRC3NkgPpNDkjjko7Ln6eIl83WH5uzlQW
5BWYRhb9u9GMUvC6XbvvpuIx0vt3lE/hg2JPDt+DVjZXd67BSzlfgmRYA5LAVLH60a/rxdlbR3r4
daRPyPvdhD1qWlv9lcFSGkhma+ZOKdCTeO0hpq17wa9umWpdE187263r9M/SzIWryfJ7OwOSGrXo
EtPpsFv+LOHemtKhiUQrggDFoio38iPvaEVBCfKA5J/aBkAIr0VAN3TfWQvx+fHZIWfO0++ox9Tp
IZ5C95jLsLvHq7YI18jVitjjaL2cIz6nLLig64xVR91PI9TsRJdvzgfdjVY5pPCV563eCxXxnB9x
CVA3GXzMytGZG+TVLsBZrKkP3vCYi7VqTI8CO7QEm6wT3rn8JRDawktoTpbR2L8KSg04UUCdH9M4
3TSM/r1iNHTOf3fbL2xohG2/P4euA6bS+oUsFUKAhkZKRhFo1jbDQ7K38dZlJ8nhtkNgM4chPefP
OWVdIfUKj+S+gNJqWT7WEbgmN4EuvgvPSj5Lf1cKCMf1inlSYJIDEeFDNXnUDzODrGb6XtOd68a0
5SGSHLWAX+0S2kPkDcEkCo8kw+qT/0ly8lITBjyQDfYJth64iz5U0LUN5oTw/f6QXwGOyoycn41l
y4GmYB9XH3gqjvseUSuCWLZcPi041zAzBezs1rhF2SgqNdsKNJCxXXmdipKPLKE00gHrcXXSLkx2
L1FK43xcGt0p76eypKNI9eUPyQ4FlrvmR8CkY0HeRvhM52X8kwDZnLFZd3EOoaDZ0xkR5GVv6pXo
l3VrlC0XWy0+fff4BYyoa0XWjF4fHT9a1nY4xnTb/24PA/giyGJa2A9R4wWv0o1ifMggGdyDrOZ8
jrrJVRwQKlQ699WdFigF837guj+8HH3d8ee6vABHlP6EE9oRHpt1i4FmnQ6Wg8vdNwqYyioP/oDy
dcFAuKJhu+44c57afXVW/2u1vG462cKonvzLYET6xAuY1yvt9q5PvibNtXJlPjPIUwqbdZBcMfF7
dCRxARffiPJ3lVUAjhUPyQbyr05yqowR0euAvqBWcOGx21QN954nNXb5L2qor+LyDs5PjnGe80r0
0aKiXsGOLkC2djqPsirZmX6M6rFRlH0D/Qso5T7yZ9YRlNRyb1T/t1p2l1jCtEn2pVFCmduYKurZ
S4IJ+2pP8AvC7wO1SV5zKZosTzgsy9K7xy6C9ArbCNd8bSzF8UKJd/wO+9XmXC/FFvquDRA+ma6U
pp+ZbL0q6tYhfa7g7ZnKoeu1vGcBWvzhCpbf4eLdDXEqchCM/gW+Dq1o/dMB3WulGQiodE2mXs1y
87wYGkZbHOJRbitqMqKhBp/Q30g5/aUNjoUlh46wW/ReOVpzOSJfGBOwFgG5wSuVjgkybuhx40AR
1zyN2ot5INThYDtUAiWK46ctcQDifCLgnQoWMioQ5VB/2iK/eABjMAcHcwieYFnwjeT0z9SIk6qU
ojsKlhd9fTBOCTCk2ZpokJqfckyD4kPRBoFHGkwgGXa7DoraRrKglfC9R0c4w7fIKplOMOy306eB
ngwRKSZiMsCgvxlne7p/mEXD/NjT85TmbexhyE2i0kCBMFQR0IovgwsSYJIWsTob7L/8bB7yv6tE
PNtbV5zVsFPG26KlJkMxgcRYr2m21ILk067kNGRELSYMjL+cpHZqjPbNFo5spwm7v82DYiz8P/hX
RYxrcBgI/hwClCQ1bLsBsiqCZoShHZExebJCRxmYHjjtWv8xa9Jx507CKk4Ag3rfLWbY1XtFuZjw
CHVny8fL2K9R7YiYglbHTGUqSPhULIUyakbVVo9xrxJXwhTcKDUCwa2aAOCD8Ic5s8DDEBCvk4Cr
dAWrONZgGIcSutv1oc3v5fTim0fHa0CxArKSZ20kCHF9FXLiJ2Wezzj7mqaSGK7uHk1zippmWsOD
xMc+BKK8AzI8ZTuURQh7wU2IetgP1qxrZJ180+8ODeT3lj25njHsz7sy2msNF9G/ijI89fburOah
a4GP1oQxR9J+ZVbL7TTVaSTZJaHtLAjFCohJMcUEB1DcXo4KQBPgvdeXpSDhAfh6VwUU33uxrbA8
O8AM3uEMV7ARfvXHw7RpkIqjhj+rNWrrX6tc/nhxCmuePepgXX0711DYEBGoK4UyWK03ewMG/9lO
UWIw/pc0fXNk1tdELYAEJwFDlOK4wgH0yDeEse6Ri/a08supDVtIfjA93/RRUpaSL6yvirSTBmDn
1jMlNgAQIM/M/rUfRxIUJ2GzBaYKPLIB5qYXOqc+pAgRADjoELQHl0vWXC7S6QAWqcaXrNBjKA7D
O+3q2P8H35Mh/UJ1CqySnXFJrJRjLn4op2Is+C7wSrpqV9xYnoDIjYG/U67n+yOJTVbPkq+1AxHi
nPGAT3zMTFm8evSSTE1VCt7v+hsOyMs4HTfAYN5J8XnuzMQscCuVoEnEvj6QTGy4sfl75cR2gFXd
LiiNugIL3hpgrx+ioiXY/iW9uDUnKsqN7DtwkspciRwz4VSFIGzV3BUr6pb12t8KKCd2K4kW81WO
waVAxXjxdlCPiEcmBSgRgo0hi6AeTNoxFz9vwfhgV9q4uQTGD61VJc01Y8MmDaaOww6FzrFbnIKz
s4hlxODEQ4Cc0zUlaZelM8P80Gxkw9T4YbbpdW/Zf0bds1jZiYRUwbFtR5R6RlGtMB2xSMYs+D1C
mtaqdVy4DUu5zZI5Spu0Mo0TlS6tW+7L+NpSIFyMRGJlf590Ws4a+PVQT9UXAbrriT9nBy7Ng9Iv
KQW9Ej7NQI12IySHTlxYwPA9d60bDe26Bp67cHLxpcOKccgD0Y+sAHDJJBY3OClOk9Nylh9ZziR0
bjz/lKzVL28NIWqQbzETifD/R8sMZ5Zi8qbz5+ia/9jn3II6jPmTJ3Ikp/E6KeVzX9aWXy8ycgx7
nErYcCgfePM/sl/y87AdFjsmSL2IaDxs7Iv5a6ntGVx0Ku2tlfq+rSQ01POkWeq9p8EGt47vXKST
zupPeV+QAbPx+iAXCTiBDWC85g/0OFrk5hOSHxWsVtRKpDyURMTNBaceCLaebboOY9iUbemcDOFz
A6KtE6Utp4r4tKIR6d4rUqfss9sYEUmrrsAfNfQxYKj70zVqShm+049q/mc8T9yrZZIs9djdRDUJ
oHliEoX9lDx4uPZRRDkCdWi4+pITmoK7s2thapK+k/554E8nZBqMie4QkMoVQ2vJjdup4mCxxVvO
xRqhKEuDVa++9/yJ7E0NMICnb1uNt6PrvOaPh4OjKw5CjKYk9FWhlTr3Cb2HH6wy+uoQbPVPG9Z+
Wrmc87vfkFsNezQ4dnMFlRUBYjt2hB7tyON0AtGtcw7teFZ5UPyVEBG8ijraUer1/VD4EKzfc94S
a9wyl0zNTf8zNciBIIb/XfBhsPM2WT4uCwTfAmym8+qCaQ0cfQkQlSF/NIQs6j3oMcw9EdlZo7CA
691TpEXCjF8aua8IV5C5/U/uIDf5tA1tafCb6N5VRBtATPAXup6Os+1Prla1fOnqwekZGVo3xp0N
S9K7/x/QFKvQ7yMTv3EVE67rhJTMwnjWhrtKzDATMJDFVhkVSzzT27La1Bu7EG0HfCk/VE9AChdM
VQsNRDf57NGJOxXHt+vgLD5wjRljpZNYDVTO86gcqvQazuqB7xIAnFfKGEaZeYnaCoO1xeLnFQdd
0Qy/2N1z86ksp/ERXpYhVcGH9KiJfykEW+ouUReVZym0MK3JeWdsagfA6yeFpMHmJufRnADm57eT
cVjBybiakyAFFRSRnsVfzF6rY9RrXvTRkWp7QFiWrfpTH6q9hu6EvQAOvnxv1tjwVZrRKkEMgNkL
bwNRQ9v0wSN6ywAlfpgtpr3+c9nWimEhWCd88K4ruQ4seV3Ooh5QEk9yFPSlV0a1pAcNidyI5h0D
+4K7HdLEjBwfts1IPRll6bfMwfUaByMOvDkYTtdNmjcuwtGzpi94bBd/o2uoD/hv+8PmFVea85ao
z1K63k9zSTNpsdg7VBcl1UAARo71lTtPJil+xd4oGM5UvcxOyEie2wpo906FPx+LSjq+f13I7XO0
gB/VvlW8hkBQDMSSvbvEGDl0eMq7JmmU7VD/pEP5cfpBoO2e0F16wntiHYXw3q8RU+o76Tex4HeQ
DNUlkN2/SSOEcend3OOmozFl2mycBZ4cfP+Ao628dczAMQrdv9dYo2MNu0Vi2A9qoGvjBPzWKUuH
/GZ8JjuGSpc7rwla/IslHJTS86rpyisvOgjH0TZyiilG+/P3c3qG1IKYmRhH22NH3PbhqRut9tDV
rzRdPN+MKCg02E/2x1pw1yaJ7MGZ6zEWfRaApDPDBTF3i1rb8FGB76cUm595tyqE4sGABsBX+fOr
srEKrAxVlUGf/aSCzpR+/wXkRUYHCEPdMzxW369EgpEF9XPyx2cjISP7vFImC1mdo/pKYemd1yTc
BpR4Vd9CsCePnJxq04PpZjNgjHyqobfGyNJWolM4ppU7XgVQG6bG51gKCvF0K6BKXkIv4wt/Rt4B
V87MSTltQYS7OqoPZUVoIi4qAEeITnFK/H4O2hYPgGFHk2BN6UsCxpu5xJQCs4uCihbhX3GqvL9z
EHB216Iy8TmLBGb2HaYZXHT1Yz/sho9Or5MsNXtAx9BgT3JsC9HQLCTD0dWK5O9txFryv9ercuJ6
CySH1p0PgG0xBANkcfvMpAQXuImE4dGp8vJ+4FoPT66RHzVKyyWI0pExVCRhyzkRSXf8Pmv9bsG3
UwpJOsb+yzpPpYp1ndc5MnoTxUU7IpKErPumMfwI5e9AYUapW0E44dqrDAc6rqAQiC5B3Ndu9GLB
BN9ummgpVZc8n1cFFrH6jwKWsIJoraSVqut+6ueRamy+8etVR2WtQlJ1nYQ5Zd9skbRbVx2ZcIr7
ApltuXfdf0FwHQDbe4O2YrgmLBTt2s0L0MrPwT+7e39FE7LUxMRLDMdayloPJzGni/Dzdi2+A/Ey
9NAynCGeSsa0fLiOs+/75BxKhxvjcGlF9Z5in/WO8KML6/fPMDDprLnGE1OdZzyqtuJoQELz9A27
ZWCQ1d6q2G0cPMep3S4I49K4F3oqTYZ6QgdlKsDzSpaio19xt34Qt3RJw67Jx0fi2c1VVcpNwKkX
wwM744vqfs0hMA7unbtZfZ7ADHgchpCikWMLsK7HjgDjKymYeH1ZhIfL+GW5xUiaBWqQPIyZ2PTS
Jl++LuYbZgUws8Ry6kcNa0XfiBITcB+j2o+9+PhdOYPyyyp7Y/N1/tuJWuwkPAroYkwG9kOPbTFm
g+/mGRV5FNeknU3v2wTDyfAImOF0oolSOj0DLzXJBqPlTJcdrQPi91eQpmN0LM0YFMeDeNqdZVdm
wQCQqVDKnIbszL78sVp1C900d0zWP5jlcZiCHa2UjQUgwxreQp5N6yphRQ5wNHElSVk17ybVZLTc
zf8JXAxP4q3Aq2W+jFBLHolbqXuP5THDkqelvN13VeaRbPUCNXHXf3yB0kWSG9nUkhYufTFyjKbL
36ieT4UmnLWvPqP4SzCuwM5Pj18VxuL61nFiLuIkV+Ps1Me6rc0TMjg2FpyfEZ/Dba9C1rSTfRNT
gvhpSUlbA7wxbyelQ/2MVWrh4cym91PcRAV+bJRtUmD3nbQ1A1VUYXpux3/GMWtQYEGw8AxxGclA
EufBiEsw2RWLq1Mp9Zgcmfsge2Kjzqi8wGdTfauNPe2EWG7Fd7iqhii1kefNT5AOUsMoiMZ33UUU
WEMuDQIlplfYSHT+6RXKcCSd6Yx/u2hu+4IyLE2BhWlc9rmAXkMxfY6yYTue8WxZNBaYP/2V+k77
JZc172UAUQ3gRwcj9n98EG/XGapJ/7RjvbJU0X4wVsv2AQeoPlA7WpyMP5+QSOJYDU+nCm3wo27x
8iMuItBkR1LuMe5DRQ5qskmRMybQrQ+iSBtSsh42sqscE01QFBICAD8YwQHTu3DbnK9D0S+463Ck
nRFWwysgyibawtKiaTIOfZHwMWn+6yAHZApJmImAlm13p3YbBct4slEt7OnMMEZoYpty8mzl7Ox2
59Q1yAd25i9BymQFHFvihyemvS7IDc16vo97boSNOrbIAn9JlDMTHdwTL8kZ7nhkjta6DWIpGxQS
5GUt4pfh3jpQdgRa7HS15ievA/XNugJXbFeuBO29tlbX469PXXt/niri8pJjjqQgCLVElR40BfPu
8QkhDsEZajn0BlVb7G5Af3uc5UfSRPJNbLyzdK5VWRUsIeSc+ltv0Wm2Yz18kc3s7RzhylQ/qu9e
32XmV57qcv7F2O70qKQFtuAyFQ9t/kBjZwR8wULayiJEGpcTymKh1TTBlOHsabbpDW+vnG+AK77J
LHuyKI9A4KXh3vKISExBLbNREGtf7xMmRXeOLCVD/s43dq7qOee/X+v+iZ81QDV3s3ANYXvU0v67
PxCZ4tUDbV3ryYhvNGVvL5UPtjsRXc9bmVk/ShcDsQQmDKy+ew+l9KpUQQT1N/4hHE2M96fXTb29
L1HwK5+/ONik4ecunOoAEnqkIX5d0eR1goVqRx6VmsEEaz+QeH/LJGu6j+xWxqVSa834FbBvgLS6
IYT/8icy/9QieNpFf8LhZwe8P+DdAmt+GNIyu8LgENb9b8o3VeEj4Am09a8/bX1QD/AaUpP6o5st
30iNtar00JzFYEJ4vtz730fs7UIjaz+eFhQwxyoiJK2S+pO+Jdr92fHFr/PXjXyZslPFnI+brD5X
kojpc2mAcGhdufZ0PI61ZuxhXpI8sFuYvuBdsWv6er/gjkqYbi+nt4BUQgyhRPQMTxPbfN+ZHg2I
ldlaR20xh6hDYDkIa7t3U2UABESHofY1VeLHTEb+zTVZLdklLkbgXtyea8JB61OKcGlQJnJY1s2Y
fn3yrQS7lreQbU3HiOI2gwmPLDmzNLTioanP/qOV+RTKduPtxI9mwCwcEmy7at7J7p1tzyJG4xkr
Py8TOJIr/Mti8MVihuBbcLYZkQNt7tKKZs5QdnkNgudW95GrC4PRkHKvss7pPvRrD+f+Od0/PQNU
dd9it3eF08Y/dTywOV47uKL5dylhRbaHB2E8XyBgiqgkdlnyCqmNS6TE6kRLi+HcPmlIyWJZ9NNN
tCM+WkTGw9IZFL52VZR5Y5nte/4Sm8m5DOR4QrPQ2fWO+3HCMldEH/y/d9JMjKwvV/HXKbompSa2
RVWXIFeoC62iw7UKZXCc8rBl2wG/rb7eLQskn7tkNchJuTe5nnFOTT6vGU48w7DmwPVH0mkSPh1w
/Gr3LgCeTh4Rl6R/oYJtDVJb++GZ3LIhXjGGys7GncHtGCHN1JXmS80D4gWHAOeVZDWS/Kkm9w76
h8lzATJ/YR3ZU70m0ZyUzECu2seT+QESiP/UJMp+rSmWec6fSUy0wAPt30IPin1zL9E9u9I4jp5e
rGP0Owz6oEvs18U+K2+Upc7GKvyLj7TzFoE6sYXSTNbkzTnmMEoeNr80o7gNp1LyaRTTWq+2Q+C9
du7RDaSKwTDsP+Ndh89ijdL8OsCg9b50geGi/LD/YY0xRv7/4RWdC0qDsmer+JsF7K0fDLplt6lA
cVzK0hoquBtHaUW1n1Vrch3hFK/1XN207SBLv1UOLmjFYOJwgK/NOy6CZTQt8Ns7SUKnY/lBerG2
x0IwTzQ06bdUUDkfFuBFHIGuwH/FMjYDKcowGvL5s64UXoAEJRyk8Xf+mnnoHl5t0jfpxcuKZJbA
QM35W2fWLFA1Zd1IKkdNpKOfHBzFYjhEXw5Uxel1F1zCKXvOpbdrFB4wY0UvexCGngqvMh2/gdlc
uKBCq2hBckMyqBKkBG2AIs2T83J0Wxa3PyUn2JjDgNxxHST40rjNqvgNRAX9t/wuO7tgKJFIMNrY
luJzR3r3r5DCxHItUqWf7zE2U7XAXDyXXUlfbw0SY7fHMVLBRb4pmzQKQjGLXFA575RLaHaTwxtj
6h88U/ndsO+WBc7gFjuZfV6PLfoOyFKKwsRG6WcNEqjaUqnbjI42cFZQUBLkYn0ilxsz3e2KWouq
txV1ABGLl2nnfdMisCdD8y35MuydxWsmWvNC9CNBDVWOZManNnTYqE6RhlR7JzbJEuXyYCEYH7vU
qXKK2w28EyrtkVPlnF+HwIjHMSDohVL3cDyzCWHcZLn5wuTdeU1p3f4+mzps0LDK7xd0WUCCnzXA
IcMcc+2UNwzPRs7qvyIA22MAHEgqurt0aqXQVZyeSvfbfyrvT+DVo8hfko8ckbnep4efz9jVM7X9
ijarB/9zw8uAd/8zmT7fKVtK5ug3+qQqjqGJh92Jj/j3V0g6XmPxp0JzZZm4iCKLuAMv/GL/6F8h
cTO+CMFUxWC/BH4L/kMRmhG3Pd+PJsxb+AeJ7im6jxHC8ekzHvc0W37gAONrFDfv/MP26xR+ZOO4
s3F1NDDgZgS1nx5y9SxtwFi4nlzmwam9RklzJSFBiYJbkh2kHG+UhcoZrZe0yG6lKx9hKPpKY4sl
EmXdlCXs1A31hIXkBEIQvKVoZA5eg8rLa/YEWgohNaQCFpId+x9xGsNK1vc8jG7CErYW3rB0+PT6
f2ue4yC3QXtd1g4m8P3kk4CJjgQHevEGs/Te9yDJ8Ka9OVAMKBlj6r2JHr1aBOCC0LlM0OUnSYXO
XTz+Uc21l1+1yJrVL7SZI2px89qEbU74XUYeq4wsrjEcGmBAIaYMas8Ln3lFxs0BmLX63FwvZqwQ
RqSDA6o7rQbAmOPOiUN0Yi4QSS+8Y//fVE7pwVQhC2+1m9I4i44qgsvBVIviMQURxANx4TqnR2H8
mB4fWlKEoMVox2y/muklDHNuw29mgJ8MBoox+gQdVEg3pafcNrUNmembPAupalZ7gD6YQsiT76NG
kmK+tuhxrLFk5w/y3fwWUv1sf4qMNexfHxtCxAMrZY//KB2zUqqZDlfHpvSIPY7heEv/TEQ4lYXV
2QhKzNG8XAiNHru9VZJLF7gvlfqsgjm/OKUxsNnwR8bVYRqOK1gesJKNX75LgnCvLIVSH3KyzzHr
XilaPHtcsb4N1KDz8+T6YalHMRLAobzOX3u2ABhIVids22zFUk+x6Sl1h4XLyP8GGnV8JFr7nBcI
5s07ktAyMyUs8P80Y9OcHSQxQF+6mT2XelxyURHYhNNKPKLFf6VUeIHmzws0HwaGwtoI4It+f92X
67LuJT3mFBTQ2CTWYDeNn/4FU5KsnED82wz56J01MC3/cqlwz6Pk7YQtbafymDI7WrN2ocgTKNKF
RgCEvHdUOSghwFBiuUJ9xk2repsphOV8TZvos5qornbDFP3ARUdaO+jB4Ma1RFhTOwpRCtPRDHFG
TXMCl+/m7grGJZqv/I/BX607Hv9gPfq2RoyPrIGwjqqHAbagXGjloKVNPdVOxDUo3yJFzqYmp4s5
qPQGwXdl+Bt8RqqcwCAr3EIbU7OoeYeq8mdQLqnQknnvMhWflIknzx5oQY0fND81cTfA2usBYIW1
xOpUMQTPtNjf9cCkRQlrrSEQgn6ol3t5LKEHhfMl9+XGNKBHk/ElrQvPf043y5QdbdNcJPBuXnuT
PbsZPaXwB/ZKeurfLjRvjfMgOmKYYxYlSJkRDqmawOC4yTF4gBeRi55+uxKE41q30ANnAixIuifv
kb+TKK1lugLJLKgozh/ghPSqw0rOz9L1jApM6LKeI7tKBAkNURrDhxnim8V5jocmfqUbovqgSUTe
TbL6jEeWyZVsNEOE1pa0exAzceOZ31esgWVjEmw9wt8hvkH52l/myyp5UCcjLAeYOvNoVgg6i8X6
Ahv6hGA6SPk98gMbbbNB6k73yIuJ6OHzKtRBDsIJ+RapbPvpLz+AuyASIY3P7bRcOJrzapg09sBd
MFXWFW4o2ymGv/ulhFq2YZq+8meJyWxMlq2+fyxxaR8zJivS2f+aqFinUg1R/J9/bVEALrxFSUR3
aTIoeE9nDByIBmIat6Z1hZUIxdiciM20PtfJQ6EfB+YprjtMsH0A8xzm+XIcQMXlc4lYVLK389Uu
Jz8P7gGvUZSUKPN9vIoTu1130nJknEcb8kjrxlIpe3maP+O8gUSwG0tmtFVAw7j0BRfZ/dXqV976
uCJsYv9vZ+O1uEioQA26dR9RML713q8hIBxlW48y7vrz9U8cF7SD1iFQg3GKO1VE+T8wZ4uJ2WsN
NRN1WIj808GUbtK26SDqlTcAW9MC9+kXKYkLg80vjsd3N0fmn4nJZ5rlG8MTeLjGgYaBCZ16UbcC
3x9XndrRS+oyeIzJ8Zwxr4IZrvJoh+dQtKDpBMLdTQclByhB4HQ7ncFzpB00z6pTBj6ayv7hx3+p
xoH13ayR5hHPMMN/jeTHr2PLik5KBI1ahotFSYaVu6+U5Xu/q+Af/D1Ce3VdvazUm3FhTMsTl/Kp
yFvN5nRbG/jB7c7vmpHfLP4iL6jcpetEYy5VG1GDfCanmyykIUiVNCp0AQqg+iNR/13Ns4qXodD0
W0Evlvb68aZPq+SKwCyD21UBf/fAI97NWapQue2GORjNWQJk5/jJ4ZG5j/mxuUGoS/qXv8hyKNVx
fGK9kWzWF34rtmKV40ZQ3aBeeBTCevpB6B7C00vY5pi0C0ETTvcSA3qkQaEC+yTL/UCkvWDZPahj
NRrlYpFrW3a4BbeY9AA23aa2r7gxPkQFtj93169SL2/KxYZwJejgZtkXx28bHfDC9brG6abMbqdQ
cK/Q1Q81KBUdnZXnexDMPeIPxhXdFztll00TVTb7AMvNGw1O8DptxR3AygPwLjzCk/Ljc6avbWkW
vVXlzuF8Wsw5hlV5jey8x5yBFTmhl2EFQMUdir7I4pF/CY2cXs7YWfZGf5W1EbqhzI5r95IHt7sw
Cw43wTNhp5iY5VjhKeOjUebLp8eDshVq9l301CZyX0DngdE7/7ULK4EWNzA3Jo4GcRHHiW1GlgJx
wpDEW5U51nk9zv6Lh3LJB8QqSCeE3xrQcP4NSqLydHZAWQdVV+44NDbDUdYDtZehZoXWmeRA4vxE
uP+PUxyJl8x8OTU6qSdL78wfLTrBBMmX8GD/7ZbsHQYxSiJ0OZv//kSHvdDOePK3n6G/XUNqawJl
1cjmAjUgQE0JBqRyPUSlZ6NFX+Qn+EPKZvTiE5mJ0iEhxs+xN8ZCReEhv15h4YJxo2xlxSGdnmzH
4/zPcQ9eW7l7ceZvyssmv7DmLytOLhYgiMHA/1Cw6Op9rwo2R2Nx04eZg2KH2xo/VUL5Q6FLTYG3
S7gIse5rRk1i6oyNpMcINXAMi2LddtS75/ZuGhl2z4467N/Jkh10LPU0hFzq439xTE9NvTVhWl1n
cbdGHbtwiU/EQIUNduolNFepvhvOneD2am11Dwc4/QRejA06tu9b/lDpJ0iNPuUIOQHyfRe7TkU4
jKF5OQdhYUuaXSzR0eUT1vzfeulQ9+rT8fRd91WdDB366UDWNsz3YMml2RdlJK2NM250vCQVTEWq
MbjL1/kxJ+TcmdSGuj+cE4DJFZypuS7NTDz2NB6egb0/EUQgwUsAJ/6h3A1tzwRg1Od+Rb7xJswT
1Wze5pH8cyGg6tKbtFtBaNQf0X4s7qWW1TZbLVFVaiARoMZ9YvoDSAD4YcCIz1JGMoMaMnH27edv
eJ/8GURHr0Vy3qe9J+wJr8dGCOkgDIsiumeldl0GxU1WMzOziYZsDxm5EX905nBPni9JKlMw3hEk
ginEu4ySShi26a2nLsxrfhFw2bmUxy7RFHrBHmYCslXUkUR/rQKJPINEL4b9/28uFBNwWVw3RA9s
r9EWzH9cefCZADM8loKHL1YPRfiJTKF37k0533k1kuofenbE3kBHXRIUoWKjOs+K8AocEcIkQ3qG
ct1R8qPeYW1PGKbV0AOiW5r5dk7tQL4CldPemoAWzS8ZaaA7AKmD4uOZKQePRW1cTJmG6gtInZlc
z3QZbr9Dcd/vm9n9LoiqVowKEdExR761nGlMUtn2E2DXGQleGAkA+BZBuReVo6OzsgoPfAKq6dVH
lrJII85DkI8bEwQyPCjCRlp1d3BOIdSjlKgMxGWymwlZ2g2ChuBp099x/0kixZzjFRUIHv/cri1D
HWn+PnLdvdvNjvHNFhJD0I69OXJUpY6uyyrxh8OffKevBBCMOESxYSJOOWcKBpnMf7bhDFGD0Wcl
SXE+umwYYNXjy6ruVZmxcOEazdJ7uXIUc3kVVBXfFev6rY433VEdXvg5hDcJXPtim7TV6uS2rcKw
RWnJKkGmRJwASu2blBsXBLZ2RXV7SUZFQJF76i8aGKtP7Ko8xdiJah6tsJxo+HZEny1GhZx757+M
uTvoXOBrOQLeoz8XpMjYBVl7KC1nGNlfi6HGqM1tx4d93LK5H8YWG3v8riY1cldmdxkdt+Esp6FM
8NbGsZfz+UyAVklIy5qwp4gGJhylsQbhF4XwtonYRf++DDOKM62nJ1qi0gl1/i35+DcCpMsBq6xH
xbf1U4jGBB65yg5QrNopU+AHbvuTF1nYW/X1rPnlgYFGpkAyQbjXgs9eIipOPFnk/YKZKncMHLad
s0qBU6XChPHQB3lbHXCA4T2ApicDwKROCU4HEBkn9UBZBjuC6HNhw5cH6V9GOTos7fOE05aHeSJv
fk3xqmns/t7u2qPd2lsHhcdX7MwdIda4vC9dmmW/ZstwieLGHFbWvoT3HHwU4FWOMSAhK3j8Il8J
t6fQTdDR576PCJDBUvPTFSFdYpkitsb/YfW+Vws84sPCMG0FGCStNCrTop9ROXoIhd3CHRu9KuPN
cFAji86Yp40gO3/RLNbb9ye2iEZ4Nc0dhHQBJd7uogL4Z7WehLxMRZsUH3rHmjXQQ0eBumDN7vC7
37Ysz5lvoukYRK8zRwjZr40+2gwm7qfgvbw1Mr+A7NBFOAFu5HGWJ4Iigv7jQ3bFCa4+px1VfscC
a4uCcwjqY+u6g0qIPPuHjqPa6sO7MJ5c5zNsjHeJLqVYpvIHTgaX9zy1LB4JaWUAuGODTBOJ4dxA
xFJsPZPyC7bmGggvaBj8GO8Qz03b0dHxkkQ6ILh9wyXK4bCEKycRUIFl/6zReX23Fm7g1ORjtQMs
dsd5BK/7vzIgE1bydxNI1WjLf58eKXEtQLn5qKzH+zD1RcGL5jY+hxdaO1LH149V0Y8n8y/9nJ2A
MXSYy/FfxjzuqTZtzxbC6TUYOhXtWKrYAU36tUHRJaAX8kSQbjMEmdgKQYJEAYOT0QcrbOPyJQ5/
FOo8EXCL3Bytv5U/bjPSdA0SN4HqoD7WE/7SYk0wwoZsGgfsXzeZcb7nbBdzrZrxeMyL15jIaTJm
Z8AQRuQmykhTF3gOvGssXwvZ0fatlKKyLcG56QiTVCPM3ggJJfncQUvidB7W88Q5Mi1TGj1tPeJq
6B6dB6oAXe6/Rb0UO8ZggDsA8NQPtqYHGWX8hQsPsPPdgHCQS7npkK42Dj2JnoG+Jk2+HGkKaUfp
C9FtpKv6a5k+0nxxH4mkZfC+HPIUcn9bl0wxi44CO9nEqasAhq3p5W1R+TSNU3kLA38f3G4qMZyw
NPSR+9uSxH/pmkdXtIIvi5q1Akh7YBfLx8OV2LMMUiywbLHq3Hk7pAGEPpf0sDAzlBUUDd7N8sTj
fMxpsOOZtD93C7o04PHZlPtJPjy5gyuaLHbsrTtLbwIE/GWHkZni31lOEOlglTJYaQHVE0dxWJNx
pxGsr8B2s7+eIiQvb+oAXpTaT5xN96/7QxLaUAsQKWw8SEsB3OOknjEEUG0goDfNtUUPZ8SHkB5D
U3WjAiaqtUwZQ+kRI2tChPPJ4bIJfEMcDDL7g35EtopDFFm1EmBjR05jOViCJPWk4GmbYBVfCeug
hOFSPVmdGMInPTLJqTSzjuy2D6/qk/NScU77Xr9Z10+Ke3No5Zzwc8pwMqvpOYERSj1eYp3L8xhF
o3qBjdM+W9+c1BnL2pYi7NFv7MLDpeg+wxZ+ZfRGsqxMco3LAHz0HPhlod3t6fd1qZOhIe6HooDo
lUlUDdSBRVS60rCfkBWC+5eweODkxuoq5ukk9nP3e8TElfF4XC4ERcoZ+ktfkcZ8wbaU6jxdKEsz
X/cn1hAErvKx7Et4youjRErfx/o9cz8nfvlKg2P/b4dgO9CkQJCGR7QpIhRmT0peKEJBh95JeWbo
GU6CLCsF/T7bxvYw3J8WeIYb9o3Qd8txvjgx+5MhU60au4AI4f4akvn2DhRFqrAY7FXTfw9C+xQ9
mrZ/iSwlbGph2d1eYsxW1BeA9oiO2AjFzJ0zi2xb8IMDa6vYsGrwMUHjQjJRHSQL1ObQrD661/S5
8paZSI1N4Gqcnfw0ZBFw5QEE6UTBcis4pJuNvCs8fDsMx/velySTrggONXAwJLe2iLChxCVkbBRS
ron9B8UmHfkOlZfNbkFPjubRqYAC6pf+567xZCIx5l519iy6427yE3qQKh2XlPHuI3ULpReWk1+3
EZw80HuO3cJ5okjK//w92k/m7qX/u5tFibkE6J19v6BAIXPXujxUv5MloC14660+TQBUZdzLmNNI
6ivTr1rUYEnMHhTXgiRA6MioA8wh/irKn8PXKntqzx1uEE5jAmvkx7hKPHOIl9tNA/SXc4Ss6ISC
ItNZP864vqPyBqnaTsK2qcGKawIlZJ1p3UklY39nYioo5rj4nMmVjFZZyyIOj/Pj54NmAF6qFfCw
BdslyKbxH+dtVSGnh/jp3qh5C9wcu0bILvyJIoBVPUIs6sOCEGR8oXCOmGAGS3a+tKOpOoi2Xs0u
ArnXN0na7n6OjRjfCBO5REZL7rzqZHIlPPjvaqvjnT/daCc+Ou8HKXAtlyp3smdTB/BdBEMJG+F7
BTP9saf/kjN9JXKMIi8m3EVeNSMtbVrAA4UzgUJCr6l01TAGzSVQiEhpGcnAbEkzgb1PI0p7wpXe
yxg0Vw4DGrJ3nZpEE15VLnh0KN/RqsdLRPh/qwaOwurLrdxCtc207ui/CfiqsDk6PWsJnLDQP9sX
yjhYa8/hldNuWF9Hi3pFpyYupLm3mq7w8kqhfrO/06LIQGO9AO6OjOISqsAKqH4KKR7MMoAq0owr
fnmlpZHWoAFNyKh7liJNkh44ADcTFhO9/48RLKgTWWzgftMfxGlUksnfvcmMXRzotABBkfEmkUkY
GShOq4F+NVJ1TJma8q/WX9mEzgJHvXXIh9Dvlz/BlpaLhx9cWqFYEEf8XqLEVS9CtPn3dSCnG9tq
Pm3EJuVa1h5xTOPA29W19W5ScKIgQ8yoBqz+a2k5yXmaktWu4tq59yKGHz/EZ7o1gqeBmP5tC5E6
t4K3og2oWl1C4uA1Vbazy27L0aPaHi5qnYDplWsAroa8KkvBr6BoN6so1BThudAotK0Ss+dyQGOE
UWJgdyUX7GBv42kywxCmCsURALT4I76sSXvFOo/sk0HTMCMQIhmUyl6nRzilpLz+wDxQYcPO86S3
uiGAeEeCNTKL1uwMwMfreWrNYg/LxLntAaO/8gnVm7fVVSqswJj3ttPenK0w7efXYizbaEdLPd3T
u2cMEnkyzJ7QcspoU92w06MfnMC4xEIk92LVaTLkcV+VOAK41SIMn94Mw4Qjgilcnb3NOk0zxzQU
oDH8SAmRjvEI8I1mJCuudW2uQmh2KO8B9y9lHjX415iYNbSz0nVR2wNFi6D8U3HRyYZ3QDwCwBZ1
krC8um9oEGo5ZvM9jA5AtZC9ANkbF6BWQhWrqvr/dR9qucE9Hk92wzKTHx+mTUftxOZ3WZqzIRac
OgwPWOza0QIl2Cw0GteY/IzjWULvu8dZX8JmLDyqZqeC9/Z36ZtvggsL96DQh1V+SUmjlIzHQG2W
UFkw5HIoYV7/GGPfj6vN+yQPQktiaKuW60VXX44o2OwQbXTc+sJ31LOk7CJFeKpLv0CJ/IvjUoTw
9150jTOTQiI1HEaTyqW4keWmyBd1pl/PWv8mf9DGcwqejVO/vn/82KutdSlUUq9EOcxEZwYdULSn
y8beMVKZDyViweJaVYuQe3hT/2hm2vAZshUSZdOEDDxtwz8617QgKdY2AiNciSVPHheC8W58Ephd
5hm4gpZXKr8S5wLK3sCuczRbAVIX728s0qgqf+BmeCBRNy+7QFISu44SH0DxV7HWklAm2jPc0GKR
oloHHaqp5BtsxlVUN6Kg+2AkFb6ggcolnhwv9z3qW0vYXzSXQ1wwtM1LnDsc8sztWobtPTQQKS6K
OTUSK68pVfIj7QET5+4IRhrTQ7/++bj20ISIJgHBkJ5XEJkvlB5vAfdeVt/pfXdzogE9UU9xWlEa
c0YBWXveQE4KbVeT95UQaUDJeEcMUrSscFbwgMs6xC3p/GcCjc6HYkCMfLJSFkmI42bF4540Zp5U
tI6lSV78XVQvqI1j5uNqsro9Exf2tMQAh4ohEj3tWGSOvkD2etcy4+fOWh6dfhNpCvH+ZioZtNrv
cMlyZYVTwhN3RXbztnFZPEKvl0rkHAt3kkpfrYz7tALDsqzyUqkns3HwYftftVOdBrBFPtpC2dF3
D+9CNNImRJNR8MQ5OkAae8gWSGFz4jcw2mfz4KuVIUpCqCoXANR128UqQH86RoGl8zimonmxDgTT
7R/lnqkHt0Jys6tsk1VDLAV5OAdbndL3gxfuR2nrGstat98JFuH9fQx5WxlCBaYBPYNy3Dc+9QBV
NtVApYGWxoG1LW6fi4+yfI3+ZeWQj3NW1MT+9uh5dM7wSOHfiRkBWUrP2eP4RCg8A8YmbHbeiDTy
QM64yLdDyuKzR1zNVvQAmRy4m4i9nlVxwMxcNpNawVSHgi7cNpdB+IGG3wUbpRqHnof+gy8cSijQ
phkGwOGdEBe0xzxQalxstvTQ41PYa2T5uum9vFB73ucAexXoX4B1HXRm6lYfHIDV6a3rwJZq1mpg
L5XUutETpEXj+e2sGD7hbC36QhFT3NIBCAqODUmKtnvLycXSvBd1EbnMfkj9hNDIJIkVYqVR0OCn
h1YXu7e6I7ukgYk1W3FiY5TDi1NlnBGiTTd9p+OatoD4u+jRCK2c5iMdrXHRnN6ZERj8PTA76gIq
h0L/gpoujedhkhvH9fMg3+Dby9eMpWUE0vCg+sAgtgNOaEQD5GwlBvAlFdgkb9deinZ0Up2wY9nc
MP35viluu7FvVYdO8WivwyzWfCtwhvVsO8qDf0vb8w346cOxIo/3mgixIsm8JNZckhUPXfidgaMU
U9jveF1K/eT1KEi4TLHqq0Uf0y7vFBeUpRj3WtnaOZfr0GpWuvnw8B2VKiDJtu7yHcE7NUbOtRsi
KnfApmTZNXmGRnXG8tByA3knd5rIBHPedZaqlCCMH8PaH0wKkxduQwvXLlccpi6hC0NkTqmzxG4J
rg5dumu6cSo8jfsYN2K6lf/jMY0tGR7G9qOcex3oZ5J86QpAVNes2P8/qpJF3zb8lJScHYUCdT6m
l+sUPTRH2yWqQJceSf7P8yX2C7hFGsyX0IGDTnI0cny8FXaRt9DDa4T6IiRAEUTRTTGY1SiOVpjY
dFkcQ2AfaLG3rg07PLEFV2Mm2DbO21mrgYD9dk5S0watj2PM9Z6iZnkrDh1Cf9hgcOW53WeeNMvu
O5gU7Zc68Hb4SLNkW0Pa1z7R0/EDoBKN7RHmfXD8JRVg1bg8hU0PdK5gEhjLtARU5T32sRqkSBqQ
tKM6tAl73LLE/rKlIfysDTKXUBJi6mmCnwuMzSIhdRZs5myAK7t1r7I+EGSksLgmI1d3LuBmx6gK
KFTwQoGR/bt13Acvt+8rw+SXq5/rfR7nnXZx/lNWXFV+HhANox/renCF1ycZRL3lONOxCiGBZmLx
qRtysX/hJV6q1h7Z9/ouiDPVFt7tGL3Z9ftBnjglqHSE7g0cc5dOPtNo49OVEj9ZwOov9br8OIKu
stnMGIwljZsaNshHSX5QcBjen98dUwTm16faQTlqSphS+dYv6t+V2k4skNr2q942onQyRWFKw1DJ
qg5qP1AtpfgcMffSi8OrE88gb1B1QHwbb9IG/EYNIl7Nf3/Kq4jx1zQz+RoXe3ii/pwoftvR19yk
XF+bY3RMSvoqQqA+dtq80N4wFyJbhLwN5TfU4yGy5BVZem6RuYooPGKt7tIsuufFQcrU1CLSjGUP
AmQ84y2TNAeqjuow7dvdpixZfo6OCUQMziwnu4k2QbCVy8nqj0EyED2Foo9zPBzuXppt/P+KZCcS
Pt2StgnOjDpm5aE7ARqVsQw3KyFfz5zL1dKrluKH59vT/Ht+LqfVtBpWPkqGwlzwSDRwoTRH9V7L
uEeNToqoMdgK3LaYCOi64wQV8tiLfJqGmwwrIA0pHx3xNJTDfbwMHswqg25X0oviY56LBXGa+e4g
gly67EOVFX4uJ/2fByH/g+W3npDUDAfqWVf6rxW9IVXFGPMe5TGdLuu1j4d9CkBgsUXma9UkfuZt
THSMpp4dkYNypVZ1Fj6vSmZ8DWjCwxjHS9YblnDILdoJ96u23iXIyIUrX1LS4sH85OPJ4BaJPmbN
U9bjFmhiZmau4WZI/6A0zjvteqqhPpblRkVbDPJYKgK87O4TUT+vr8TcACZJ33Be4m+uzgep5ANf
E/KXPhot4bFuqrxkhJlWipHuD0+K/K5BhLTWYMe3radvlFprS893Xn6XbQKpulIY51VLgd2K6CB8
I29P8M1ijrt+BECWF9f3yT1rAOlhd2g+ZnkbvPLjrIKKoif+koqQ4Opm5JSQjAwJpSO/iaT6e1dP
/uz/IPBUJ1gQuxP8D7/95m9Z6F6CkDOe5QlSAFz/ufXpsvlza2KNxZYadJyDq745hr+uLWIOvXg6
c/JlgdfToUkM/y5+84830VUSBWgEi5BTPTgloi8bOV3NIWuhq8RVWrirHQjn9kV6iHXdvpBnecDo
T/d0Y0zFnpk3vkgoQp/GD39LAqDVNBkHfQzYotQTVkJb74VKs5gz4M84G2StY2Gs8BOlDTrdwjx0
v3cfe2UnH597Aw5eXaBQzMiX/E+XYu5CfI50ToNinBP3OU9ic77I+YIKnVle7FmI76ejqqraOKNf
PXCT4ldZsVwAudhoNVpOYrBk3oS/Mhvb/jzeLTQL0uCmlgI/lTv7oY1toWUldRnM2IOthwOMLqaD
3fHZRJ+9baG0tmd7QZCO0XtPw2a52eEBln7r5idaBlRrBHGhNIAGmiHs729zQFRYTwclpnCvPSgv
zm3wH7nv+UhJ7zcslKdIS5EpBDubfVCI/QLsZnUkQoFR9Pu04fGIL4k+a2PXFAAicLQEEITca7NK
mdkz/m000Bojt1BTZJB+1EPtd/LacV5LkfSSZhqS/7923CLIiZ5s214gi8B3R5GbUSfVZ0Rqoq56
H7JNzvGRC9x2gtkAXMvUGM3gOi75DePy0ZYAHswr3YK6pS51NjVWKxXzM617tDVjhnjC0lxFzttS
MkQbHt2ZVprQD42qNnEPXF0mH6MA5jErW8/IFOxxHjUfop74UigCtqUoaTy7YWogXXKlqNemaLsE
TO2xHACFbV9bjRfwt1qIJyrNeO/3FIZ+PUwrjpj4rRPtunmBYrR22lq4yQ2DURuWxzyKOX/V6F10
+c3IzJz7rA+oFyoL50FwcTmcO+8k6vbthYmc4xvbn8lxs8aj+siZ4C0ibSTt8neJ7WHRZJ6ve1x3
1bxRDVswp6S2klrVCzNVizTJmndVCGbGxSz6hyZQgaruCsKCJVIGomc2tUh3RPSYdZYRyzTbSCeG
UHK5HoRShigwfo0bK/TTNGge9e2jxEo6k7LvHEIK6iCPXlWPJrAxOkZV+mqW5fqz2S0E1Hd9S7Ly
BQ/PqRwDwjuBPuSqCvPx65koHcK66tAEbnfLKTd5ZxnCSzBYC5RpbtyRsjasxNyFh7o75DoRIZ75
FYme8kzRHf+B6ON5qAzqBn0oayc87JZUPiK9B7g/JDZJOPWhc53++yapzSO6THVLN/FTjbeQP/WO
g9Qwiq4EYtSSbXFMQtjLgvgWiR28aeXTyocdVwutFctx3qpF5EDTEDT4P5L3ltemtLWR6Mb+eUqG
PcXXtvGyjbsn1Gt/Mq1bqYNacUwCOYXioGfrA+GIdetWcrS115E+ID49bHFpDDM8eWImMO3CEkvm
EwNsb/teVzTdZk/6vPdcP0XiH2SAFcMVZf2gJTGkwOSWYx0fiSCO2+OdJXoREPftwEr9x6wQwOch
u4seR5OOvbAmgN8+VSyIy5L+JECELRPV0BtzYeacT4s11780uKLn4px60VtToyXy2E3D+9xrt1Ya
OK+I0QdjBluWxMfvqenvlndpOLVfpvV4emhwYa9QtZAX7ukcB8W8J9VJ9/Shk66ggwuBhFWtrTob
C45H6pnai7cq5RIMZmSd/ULMuhb3jMZ/yMwFTKWBI6pJqSBoS9a4l/m+k2ovnVbi5xm+kdofnrkp
wAARHCVpvVfwylrkHQ2PfJoXogNmuHzDCl+LMNutMXL4g9dt5uPzETlRvABCTgI2Vb4yL1JluFJC
YRncbV3BREK3oMnaYDFkHLPPhF2PMoejEUp52mBQdh5feMCAKsi/FUO9OAVEDW0sTxrEhPkmXP+Y
/oGHIlynBzdmUQhpJVlMp0I+WVxOT8DM7PFysbjxIHkl5N8YNcGlqiWAoHtkNQKvutHmGaKFmtGt
5ZyF9HywjlE5+9v1/cQMeAJsGG7YgpyT6LG+OcNogyHbpIVrI8TNZh+oyWyL5LfJ62nMIYrGSz7G
hfmHuFv2sYOvuYV6BuV5Cc12I6izFFmPud+UqZUEAZbTkOlP9JPqsuihYSYmIVN2BMMbW+aPQ1n3
AZGlBgnEA+JZNKJW6EkAmmt0/jzKphqdj+VNZmbcCApWbokRCj/vmf4DoPZmS/6meEzukOGWj/pd
/w8Leuxg0N8RbtxIf6R1Q3QGnaRJBhz13H4PVQJUUfTjuMILtfrpWjtknzFZMk0w1rzqdl6MaNKp
v6CdJ3PMEN5lKZUI5yXrkIs93apWEoYWO9veutdjMsWYt4LZnh+bwAJpj9TorptzmXEn4gWCteJb
T+6SqBrf6CE5iHe50FrJ9y+ALSrm6tzAi1EAjYwhQhSL06WryTiap2eRysziCA/6lt3dC0V7/ELe
KyitPtMkmgnKFbLwmwH5kf2yZTsLXAW2bvNCMD+nOgwF4cpO55E2/+A0HaRw5nFmh0xOoHVO7ysC
HsY60y1iEyx3HvId+z5uwKKLr5tCnxYvFmArPcROKiPj9NiIXNBXw2hAXS5zg1sqs4ZwiGiF2An5
3x0rX7+lYWaf9JvZzakZSbUPz6J65HAI6UMxXftRciN+oIAPUl1bOiViU0GjPR+wD6n75QK1olpG
7zKwdXDlSfddfSZ0Di/LCSzPFtQqjnDWt0Fx+qgnAJXqe/p6WBueAWc0la27i/d8Bn4KaXU5mldQ
OAe7B+F2RXuKm+c4fZJqCGJLYltbuVI4JQSlk/uWtNvmyRwY7Wvk/vG2c0blgaXSE1E9gstA3ml/
V8ipbCAwXbxR+J+eJfqaP65dXpWW+YYy3VkMgQhv+0bbRma9q2HtIOTIiRYY1YqYoJahISdoQBfS
H9DE2u2Z7IvXkil8fwz5yC6D5o0IkktMOoPl6AVnXuKm79lzcXNKPboBuSVI3G1X/9E377/hFJkK
rahJD6Uf7uJyJ9uTf/IJSc6NoFxw4YieJs5Be1UcI0WU5J4STc0VnCgdLVIIHDXIAr26AD0VmamS
XZoXecqhDb7OY1ohyc4eT7p8HSpyer+biL48B8vzqwB8OZ/0QwBbISQTsYHOEYNTXPH8m9WsZ2J1
b39O1t336XIRHI+z2BFjphyvJ/z2rca1YmvV3FBR1qTf2RqZLZy4AH/2s5lzHGdrdkBLoCkSOxd1
M1G6RDWRhvVZxG/ehigxn0VWy+YSkB+52pl11PjnhmYtkI1uBqBiTgJeC7KwXCbWZQdlYVeXgvr9
SdbzdEr7T/XTi/SAWvq33Ld+aHx6SqpnCyWWw5184H8FWwdr24CJ6ZCh16bHxQoDXYV2TNDoL7Xl
ovvzJ8uuks6ut+ktuicJLssUHh1DMzoa6mqAf7KvrjGcKogGtPj3QdBBsGHFn0ERSCm0qNJIJU4e
nSHoBcx/nVHp8Gr/zL3UxVOVtTWeE7BPjyMIizmrsXcn5J6botEca82jWb7993wWi4Dz11Tb38MJ
8y+LlDMP7Ul1KLl1A97cuvKYHlYSdHnpV6aulMdMxOPmg1tvW+mOum0747VHCKZL3RQ3eJszLvsu
xxoJAt/Ge3J92C+b+7zIwUP29P8HjmdYfuA69vwLw3qyTT85EJcIrsNJidFI3Pl0ZquP6zfEoOxO
3GwJjGZRj2cX5Cw4TS07NMqOsjS56/Ag7h2IVSzPYIgLpr+B+pgm2ej1reM1r5LgVMVzMuvHxzW1
5BU64uJauUvJyzn/bU8KTKxaUnofoNyR/DydDThH6gO4E+82eZzMmazkW1uuwaZVse/u2QugHhgA
x8CfCy5PlMIjJP03c5WKyXQz5yGV4qS6lth65KvxKt2Hcm7eI1fnJxEaodKo/ceTmSGQ8RcEwyMi
Lp3xhbppbBIWqPMOOCYD3BB+7BMtcXsjgFyKT20Tit9CWUi74zZ1ebEVEAIM2Lt7hGzzqo5dIM9j
qBiGE28ib66mz2tmqTHmFsClG0w1ivaTgyIMB43fB4YS3/TO7xhfNDskexbqv6Uu9GjwMR9jZ43L
FvCPTQfZ3pHtl5wyjc2HlTpNly3x05WNoS4D4vSzjVyahPl7WNZgeCyzU+qWSVctzRPkWnW/an8r
fv3VUirIh5qvgtWqwCeIj5lpwZe+hfknj9OSN6a9mAuMdWOmJhGj2PjbEC3fSg8S31V1Vt02lXlY
hWIVcGgUsyo1+0hK4vXTVxAK9/fMuiAxMngvB0/9+CR2lnv2RDc7meJScJRmtzYvDGiid1mpYcgI
EtkCbSxyKWVwLy+PhscBnBiRCFOZ6jdqJ16CtBX54s0ymi1IWVfl5W4LCBwulDZAVcT2VzuJa9eZ
Jt13/EQqS22Ru8thRT8Yy1RXQqRCoOHha4OYyQpAARqpgAcG9P2Wh/hF47YtqNZk5Drw2JVK17PN
9iHCUMVIzPXxoEuVOODqYcLHranvvpRrSZep4BXT3TtdgcE6nBsJvVdmUXoxSDcxrJ8HiZXIGY2l
VtQ2wr9aZYypjmszvsXZgDTKuz0S1JQV8gg8nd3fLBKnxJgUtrV0WYU198nkqkdxiwXrQdoVEkaY
EtxJi0L4vO1gkYM7RfJDFkEodAY303FDNl9kztSn04mjajYZpVBwiJ/hYclSjx3Y1PTF2IuxVNxn
O09TPCWJVSc9p21XME9Dh2IHXR7iPKgsfE1XbekQmKLYs2hht8N10IscsVVlofu8KneQxRT1tlwa
rTDQa5x2s9yOu0c3CAXdbls0JTsrWPrT8x2t+rH6B9ZoVJAoGVpgJ0iQKJhFs4DiE9AFKu+hhxQ0
c+KxU4hKs36hZFqjzhBdFhLGwEL8yyz0YkVmKN+g1EjrOeHWx+d+viHCM9Yp68PprX8A0WrhmK4I
9+gPvmWFsj9dnyf+lleCqOMdXLuQNj/yp1OXn2IyFE+yJtNadu6FQPfwf134z3oeZr4AyDMX+X/s
ub5EwjFl/tIi6nWrzxfnjcnNl+SRIOI9NkIsIdbDbW7EJWwjMncNRUDUiipZdY+UnkyABSaJaSSU
PJScjvpFoOtBpkakFlg3M9T5O+S4cNz01zPYsvVwvb0cO2zTkQOrF28p6mtus/446FTSMSZ92ObD
brDc3i+uczro6K9L3fq9N1NVip33FxfhHiJuxCbgRugjne5Foh4XT920yHi3UswHF9UF4kLjTHu+
Wejxl9qBTXWKx9BC+dqn3NK2cU1t0LWFQagCyTb5IhM724HEoE4w6TiRRlU9oWttZNc6PUjRqgdP
U1V960ackTHR52RVGoxbBE95vCkeyPEfkHE3/4qgeyEM61eZjyO9ZBaq//UBZZZTQYfVCTyPirsj
9D8kEQxszq7bUCrXVhYmx8v7tFXQKG9qi4NiLIWWZy1eHNutwOdIwu9bmBI/kQQWdohXphCxNwyW
blLQZpEj8NmZzoqXHEKqvCwe4AEgZzDp3eQAF52GCbw3WNSeW+oFFmGOwPOG8SH13CScj9M24+to
7tMMWaqFAMbD4vRWG/3eeHmm0RLdpNuOnaY/CY2mVVUKU8sAcuYaoy5vhCejAvfdcUs/PI5HSiLm
WHMAIYCuKBcd+2ZSwaCh2fud8Z5z8cnb82LAYElSc8krjJrqGchkR1ZzXSIN6eUAmBes+clqe7lV
CE+AmTHE2NPNpWxwf668JcHIHWhqqDFcVtzgY/EKahBvxXyIuVb5EyjiJczxLofaa5r148TdrJJi
/DBgojbUx4caCZotB1SMEDJDKBxkE4LzGe3X3/d0tnjqU2f1J9Vyb8gtsH96J9juW9SD8aF20Ftm
dprWIL874ojb1c61pPf3hmiAS+3tX586kd8mMFYGOfmtjPXUaoL0UGSpXO7xHF0++Jh9KXBMdHrb
/TT7m2wSSrJenaSoH3nKYwRM/GfdL8sNVr1g32JoiFDPJrcghomQZ4k7OoV26jKEMxDTG2eFjnhM
+vbYXPBqjjdatgsxYuxmUHs0biqEUf6SXbElW5CRYzdsVk4IjFac39nPF6n0q/N6EXOknoJYqPvj
vYXoUzCmhyn9NLi32ZGmBd3PnXIHxTJXB4a7dHR+PxbOcUDCQbOlraFYVJJlPUFJ8iegK7g0NGO5
MuZyLLjHfH1PBgxjHUMl+OVYgKmBTx+xxHKJrfeIio0eXowEEh6XoShh6e3va7CGvzPidm1WzUIo
jOABEsErAdoc9twLfUFEeZvG6OhhRmrTke6isXfE/3IQDMo3WQk9rHXwXVDG4nUkuT2vWRY119V9
HhNEBCBWx0FUbtYl9ik2RpbbDSGfexdW/7Gmxpi3TqYaej/v8kPoR0z8uWywwyNmlbDvt6wpoo/G
46AOt3NQ2fOx6sRosayM/A2bGaqvFSStQJgxJy2ji4aRj/4XLv0WcY+JXGSP8H7sRMHoyQ3osd+X
VgJaXyhxFeclVENK2+YwNvzJ7RckNsc7SNoA3raJW8SXu2rRMIO5HRi4bTYV7qWWIUFh/ml1HUHk
MGqr9qOzCJRtzsKqz3TuH5m6cXr6S5h2WfuWthlDhsgLXGNu3324Hs72x7JmhkrJe0GXTTUlgE7e
8zDvJQZVa2n/zMGJZmnXn3Qk3GaWUx5kKDGCAeUoksItt+LlbCLHbewc2PtcIRTnHvXuqCLcmrca
sKzacWZhN8R5F9tWMXDAR1NILiWPIzynhFdNPjzqcCe+nAqIOoi2Tz43Ks/WQQC71MSHG5lvZnUl
9yJgQR/3ouDFRv9igZJTeUraUXr7cbmGy/+RdhxoglxC/drk+L2lysnFHp2jhJ5DpgImq5Cc08Vs
gAm4tdm1uZuKzuzJU4Xgk0WCr1gXn215EYUB9bAdFSl8Ixev7klmaYxU2w/v7ImQ8AUSwBHCIyIE
5cN19RJoTVReaY9Z/mYJ9hC7onCbJgq3PPKDGLshy7p4KtmAl93HRc9fSuimu3xfR9I4NG8GHsq3
pwyjlPWR9ESrCoxYFk5LEQIbNX0cx6c4UzMjNNTVj335KNldLZ7XCRLCpv8iEkjghJmepNUweRIv
vEaFDIuZJ+ormzINcoKVv2NWSdeS/B4ns6uO4+1TKCSiyjEQ9muOaL1cxO/KnWEKunNL+elylIeh
7YT5+NQx8ak21vMNF3V3VPw594zYu+bWAhhSqVimYCUa2wv65Ti5rqJF0lBaegABUkgHkkSAbrkj
ed3ahgbV+oA39Rz/Kqo4xueChbMMyqAI8ng4O9zKEzN4qohjyUKjIjNGTFImkIZDackLLAgbj+B6
6k5GuQPZWC+/REKPEOTqh2Bppxl4G4U3n116ASjGSz0jDxbPMkumcA8/AWp6gXy4QeYo7b81FVVJ
PK+0gPXw+pt9g/P2p/eEdpP26FuPClMFGLJ9J0iRjrm0ZHzNoUHSVpIjPxamcyfK8H9wZ3O47AWc
H6u2UJPsJdg3WWCTqXbD0eU3ExiTh4mdKxI4aDgz0+yNY7ZOgwOvOF2r4BhyCd+p/j9dGtMGL2Yy
rS5EtSFLLMukfrtBg7E3y4x7RElFXDAuh77h/3sE+sTmjRES3VK3+mCzJldioxbJJBKV4PRcqDHP
dyvGNju1aEztzUE7rmdoafvKRGvzS2YGr80v6dqyDVoYSCyjmld/Rm+FdBHbocopY2Byu/GOPlQd
wPnI5v98JjCkKJ45lhqNwodTwkpmUYoJ+KWnB5NyWifrUeQxAuyjhYQ/Tx5Uaq+SGIbdH0G6k1XM
s1OAK8c76wkXn8tWQ46CcD9TSmH5k4LxWDIyPxKyL8B6/AGopi2sks5tC8INNux9r3i84Q1kYnmS
AA+05ixDiaR4Kfj4usQvCfgbjuz1uFMGxDG0yKu9hGGLOLteo0c2vCVOGTXuSDeb+ollwWU71fXl
PjVznOnbB5fY0kcNwxji9EKEFFQTqaLx0oyify1Lvg2MjY09Ph/DcwLIOOTgsKlEOuWjo1PuPYdB
d6PoEi3JQ6GJmJRZWZhWR3e3e9DZwGgtRORBh6Y71UhDZQNFZ89xBerW6v1V7zTMNzo+4YsJPjYH
MVGmLyi/JssZ5SWvj+MAUTVoD/quwlIFVX+v5z+2yyxu1c+a0Qw4INzDiwkv2sF0tMWt27beL41J
JKC+6ym0E2uW43rvmbVW7+bfesyJ9+u+yN9yF3isvVJASOYYwIj00RYTQ37ur9sFS1sGTHRRFnhq
hHBNySmS3gNXe6nEePwsaFyKtzYoVQEqjLrRjW3D4HvZFKe0g0Qb9hTuvXNDAqcAN9zDZEGgKzhe
0g2/AKS0zuIKuu+U8NYC2w2ezV4WvF8E7Mv4iw9phJv5/JtWLEpNBhXIz8jbs0Ke4sL7QlvcWjXW
XAxCU49uKLEbh8vlwNNRxF2Q6AZIahp7jmi58IuzMiSsfoRAPyAWY8OcLBCrofdtvmx+a1AuzMOP
ATGQoNGrDqHHBdO28/kdmEWe4r1ks21JXF5wmLypla9uzBRHSMkBKboMeRj4lCGAvj2CN/7jXvS/
pW9fXOXVQlkPfOOpuB04BHhqS9HJAmp5F9OJUhHr5JIvcH4gWwSa62XpxtJ8GiipS7toSQv8+bWQ
1CCUVOh9FYP7YYP78OLfApAPJaTPvN0dVQ94wZasD900tygHUY6oCIbBSNNrYX7srEpiGgwvcXg3
6JZBLgBSzLa+4w2Q+qZHMvH7YC+0fyJiFSb7RqrlBmf4PMXxjsioXrtM2wMX1MteZECQQU7/qHWo
D7xV//l4gFkXExHalIyJd9HVXRyRKzlJ3l2mkGaVQzwQ1ZkPo1vKQ692m4mN5qltjuUj6p1fnfvF
4AbC+CHCrW6Fccom7thPBJb5j9OWpuRe2UJ75MaaZosnVoaJfTlPZEzX3TXwovTSxXJ5YnQbGkG5
HOSKq+H3kP0FtwVHF+Zs/lm4XwE35mKZDXnLCD4mHhjpvxpvA+3WPLd2Z70rIausMbwve+sNFVaI
LwAsDFH/6ingS3IrA79GFDJuJM8QT6eHZ0xAlHLhsRV8mCYG0wvXJ1ii6WHU9xzJY2BlalgdADlw
6d2/7cqESXix13CYIkF2mrcG8Xn9/NuUvJzA9wkr6nem8h8VlQqnPWZoW0Uw5vbelp20K9SUFhKw
9Akm2R/0k/YRdue02vViAJoVRCfPkGGRyJxEnuVWRyCorXq2pHbYGOU4dLsyBQuxhKonwnSC4CEh
D3zecmv70CL8UQjgtJ8uWJLQsLnd5b6OT6+plzc=
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
ga7z3iGMhGhga7TzPGleypVOHJn9S7KEP16RJ6j/y4QGRddc7/SJdXJ2zPvm8FTCqWlJhu6/s34X
gPP3kw7dN1YdiZ3wZ0Vzt8uhC/B62KTkMGylsJT3Hm/4AVsby+VuOus10FHgOgp78G6FqJDW2hD4
FEF7AvpJ8kF9S1ZR/yBaB9R5/vEzgMTG6H0b1hzTpBGPyaW1S33KG60mDs4uY1wSc9WkIOuDsX13
gE5v3E3AdV0s35W8mk90srPFan8A4v9WhQvKv0pRdTPwajKYNoHYw9l0a0ijfdCCo0SwbSJr+KOr
7KJQNnQdeGn2Y8dg3BGFPO1H0k02bZuSqUQ8rQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
dBwrqXpaPIvc4b2fzIcAYNKycDBKm/hw0N9OirP+O5J0w47WHpIJLrz+YZdtlXZ+W2OT1CCdKga8
l9q6LpHNXfMJe0tSBaUQJS9kx12QCBYd7pz6Zz4XteULmwejqAW/r/1SNtjKdsFfgoOhPbvsYv0n
RR9WE79+rnvNSo03sWloLz3If8EsTQUj+4AuHA6W5eeLCFFrjEJDELred9ftNf+GjbKQ4DD9VT1l
GYpqKI157tMW7VzaYctB1tIYsZm6N1scQY5/pen6aJE9XG/GVJc/lUhiKfjKkAB4R0V1b6xO6o/L
Z0CvpttfY2ekIVc0VuCKq5gMTfn8BkW7RjZNRA==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=9072)
`pragma protect data_block
3MLlIGXYAu+SNVZUrN9axPWxB76fSavWP25CyQigoZQ3T579rH2tX4mOroKAFnY6MCrE4zy5SoFT
o9pFhWobhy1JNncmCcy/a0fRL9ZlIyjwjHAt323ZL0R5G1zw5cvTmFWPoZX0yo775l85Oj07XBYY
i+0FcCRCKdgsQGwhMUnpc6ET4ttBmjQUuxB6g1Afy5ISJRNYs77D5E8aOFrmzUzDFsE9BGcX8wUT
bT4zFmjkBZBQ+KrbdhaUiVbninMVuzKJe0egFOCGcc6CdMPwZP2SxWGkscRsjPCAUdXGIydg5Z31
50m/zUoKITRK4jViYvnHt4f6sELIUTWEwPvxSg4M+j+wpDH8hMQC98bpm495w9Lz7AbFBmLBe5IG
17+sbfU7k0MY2fUrDvsniZvkyXNkbKvNrkm2E9MAmf3uKtqsnMU/tF2um9tYyMuoXrnv+cf1WHME
rcGa/NDEnGr3zL8P+jWgeThli88TgswwgsRldtZSZHdEDO1R1Eb97kPR2KAaazYlo2Q2STr+5F6V
SY1q0ie4TtY/nmeVptSZJNGauW3hhgmAK4fuCh0LfgbkBsnHNuCX8t9sRAwVUkoEOlvg+hIeL3ch
IbMuCTBsi9ym1EZ2NwdIt6YMzhAa6xgt6mL0uQSzppyrK9CSimYyzPbah+kviBaNcZ+XJClYLFwg
Dt034rBFaffea3MI9/T6EckVHZwmBgwvpnfxe5dIdxVZcMCrn14d+8gHoeJtodrk7RCejHv+C9Jn
yRjIaiu6w3mbAeAL4r66PbCB+S92jMdnwdBtSBcwI+pRfl8Y1ZjnMUax1D4+e4G/2vS04zWOHJPK
TAm5M/l7TRLujzCl4M5tq+MN/Sl/TrmT6Z4/ZBXtoFpOHicvprtU+bB6bA/TDiQ+wyauUCUWMDnD
F2sWssLTcUSqWyGH8nZQJkJU1GRznsjpDp4OUZFEoGr1SIfqUXOeUdRWE7kTsTGtuLLkFRULD9ZC
icKwOzgQXLWvy1haIHsyX6SZ+d2z16A+qjc4h9yGuTAjU8NLa0V/nk/gnsMB1qd073hph6QLxLJK
r4sFXdYNYgCk5RaS44kcalofpqStJQULijgevhq0IIAiHku9ZgDSCzWAw3Mr5M2bNizLX2XXA2zw
yD5SKKgh8NLJ62Z1MJq1d/+XEurLezROXf2MzGpmtx5eT+YNTMToyw4wlcI7tOteLNTVwpN45tUQ
B+wyQRROLfJbya1slSCz3CBx0TkfIQfh2iiO78hl2uIlnw7hygM5cDhSSbRATA0xa7ahqhvOPN7M
cHlx2JtFdxdsqSaZD9QoJ639DDyU3Hou+ECwMn0csUSwgAS8rtGVdP0Of14CplgwrGPXstO6akKA
3u+imfQ/w8L/PLKXBmZ4JDbURy7k1H6RKbw37csxd/ZvrS/pSmIkcNCzp/c2DuOoQ7gmrvF/T6P6
o66nwV4BSbtkXVm1Gd6pj8kuzFas4d8qUgIJYtO74n7f/EHBC4KRyKr547xiGiwhk9b9qd0mjPKY
rhYsYy9gXuZh3r68RGneNEq01MvW6g9QFwK1ZOIvZDYOR4QWzSf3jaria7TfeR04B0hTDmN2pnIe
G0GNQyny7szBaDLk+3oC5dKi2x7IBMiFePNumBGpRQwF3BZOBafJAtsThr6J0+IuaIyGTu6q0CRE
pK6/stbZUIyDHLZTtsEiDvCUoqJt1Nwycg1jZabyqczbNym1H0NA+utNZBXESxVE+E0tL5xp64UF
6UUd+qxyLwKovERkzivDR8GuW1zTirEOV5S4VxepjAekJHQRl/DLLebsO05p1WmBlr64t8l3I2Z4
eBoTyoAckywhyY3Hef2UK2jwBO8dnRLD1Fu46o95g5M70RM/CdS1OdLKSF5ccJEDtzouHFkJV1Uj
jF3ui454vNAg2ROOQ3kKuyo5BsEY2EVCu3TpZq4c/q9GQLsRGPOnx3VcTR+6BZb9QBmDwr5qk+/F
Mfy0nKqqzp3OK73AWybRMjmJczTm6ffP4zxEkfUdzR127EO+OljvRItBn8LSuKgqUpIu2NxDCg+f
A8xmKgcdP5Vj8cz+tus1NipaLcnS3rd6rslS/DaabQM/fOpx4ERbftZUSiDhPxRfGlVjhYH1zMEk
pr486KmY6LfVGaqc2pCdgIkuSoohsNiPN8xmmK5O9HjxRm7IYdaUIvotow0YeYsJys+80/gJB5s6
cE/ss5YkBWNMAqtri10qAqP/lHRchjbTFTFInn1auRmyFcN5WTjU9MqXhbmBIpJrVs6hQ8bjrGbe
udyynSp5mkE0eE/e2v5I1wi1YhxlXU/wpSQkq7AW/DgOKirxvaKomORblPuNuqND5ETjQo+jpEPM
80/aOZIyPqN0aWmrTJE0jsjxS1AJ4MOENCzTG523Wq1bgye8XzrN4fo53VpdHD6EPKSh7ZgGV7sq
giQ8mzKHA5CetG2XXI6zrPk7Oe4z8m90oe+OF3HP34C4sTOp/x3Y+GqefIC7NoHPNtvs6PK4n21W
QJDfypWh5VF59VtNEgflzAT2wYDVtih7VEgDNBwrj5ychDhaeRx4+0dTJ9BZTa/Q0qZqOY4erpsq
jvneKxGNPh7zRngog7RWOBuH1Hi9ahuIiY+gEC8RxoTw0q9WCloHfF6cK42Bey41W7Nkg8Ic3W6O
AV81HlRcI218/r7yKU/7urKe8KAq0lmfWI0uIobow6NRr57vlBBhnMIl/DXynMAD0MicHsH1Dhyn
h+XWBoQuDUWkaHIh4zZ/+1qRMEs0NnSiSUJpOxoccGc+tyhoKIypXhHvUevk4IqtTmdXqAG9BJVV
k5OY9fhhlE2OW/ibdkZv1N8TAqzbACTxaJsG4yd9IXNrWQH3memdIJYipNklf5EjC/KvbTm5tyl+
BLxlplNCoR4T5q2klsjPNTl8nKAiMYCZJ29rISm9ghJjvtpxxC7iQxNuwy8DpjfL8Uf4MMBxii/H
GSJtEZy1R7DGqeOvCIAWAjS1+kkxdMrlh0x3ruEo2+mWagYuF7zcRwv3TrcxsdpZpxjAK3KuJQ5d
X94lkof9p94Q9FjBqgLyhEjFTPbeSIdMHrEiuPoqCq/SHstw6UAe/HyD6+3m2O2WR1U2m9uPatvm
sJxRvmVVaHWurvpn1JNRY5/mpZqXlkjzuf/rk4eL7YaveH1F0WX+Ql3Pd0MA4RpPOCPoYJ6ooi3X
oVoBCaBgNLwuE9nJoaTWldtbdFa4ZaDZk7rQMlAKVWXu5XPEChTjxfzXr9iZw8Qdf1rTNBPLxMWO
LS48BLsmr5GXjy67UEUXHgGbVRrUX2AYtWS9hX1O9CEOcvgQiFyWG7+HS9TBB6SQ2461BLLzDSIm
tHQ82QNlJVtLqGTo0WcNrWtZBNk8qWHaU3vXA5QOlhzZmHw9E/y6jLn511lV/OUgJnhM+VkJUv5u
1GWSh+SGQ7IGzBlp1mAMXXSKsY9cSzVqiU7ytCkCfz7j3DJH5ntdAicnI7krHr+QdHoHVl3cPRNN
NTik7Oj2TIhkPWTVsDBGPqiRUwIeX6/EI9jZpwpEEOFrirGLMXLQlE4bDVag+ARha7L0G1Qn/UwS
ejMGqfZQRAgKydtDRMPe5ZVBcXjxlbFRxDPhda1EEu9YwjoxssFUFYaTKNMkzgd/ILMYuoWISXaK
+L64nS9GUjgI6nDexUaG+DxiNSa9V3et6jDkOQxxrgWcmQBpkk37KtycdmM0jrStFP5wmOsnlJFp
SCGPeuT7Jqp7MdnYaR5o3vKVglmGTbwjVEyEhlWMC2Bbyue7NnT/dyA0LgjQbOF69e2BR2bdmIIP
aBoT0VEoRqavKJW4VVJaM54H1gcMOvTiiwzgnJDFqLa7/UA/7wMiCGu4uBnB3/kQzacm2hlKuJQf
T0+vWNMiVBUy2cr3ft0/kuEG36VBq+hWxfKK49u9O1qhxvIIn1z1ZWZZD3MHuAZXojeGQbtv3kru
U3XT+pJVLh5oW7JXXxSWdaz2//oEhs7UgNjE6GxBsIMlGPBbkJ/ycx5yfyxee/gm59BlN6y3qJxe
INbnePJ8joraeLI54HYhmuIWx90XFHYoDJPGQspHtIFbLkbuwDmzVGbD7LA5GRjFnNUrTZfAP1EV
adRX/fDuSPpw1emPPqmQZH5VK30d64GZveWzK9i1yfrdv5e65TEzX6LlxttTYQKkEP+dtczwig//
R1YueNMWN0TwjToe2drBo7oIH3dvjjmCJGzj7L0KVXsa9T9OWhDmY3bFcKwLDrLfrOm4R/IuFEHK
WOdLDSei1hDzy7wy/K8jki8xgNIqCnChyI0UL0h7MGpoJZmBKzpmB21NrbYCdS+XnclyZ4pPkj97
Ylxo6BmW16US+sj65NAvt7uBNJHj+3T8wr3qBqSrSQsvZLNHSB5/u+5ZrPQSNqbhhjQv0NxUm8rW
8mlir3nvxXFJPZ3K+S6GI2Qwnf2OY2Rw6oMPtCsWx/sQiTfPQtb0pb9mnbOcVNeiEbHXgFZ0MLGz
HSxuKW1kexbxYUG3eu6vL1dlUHRKIQ/2irLYTwymVewOAwSODl+75/uB8Wo0kVVvpXGw/mTINAYu
7qVxHRYXpj/ksW4pfMUjP/9kM80OPdcSc/1g9yUPA2RX7QkGwH4JCwwFsIgv1mvu601jFz0O9Bkl
0PpkocFdGAcJZC9DhmjGWZD2cCN9j8QnvkQzeLUERyt2rqFfavwGkaLpxkfrv6OpLM+hpop9o/W7
f/p/JrT5qiANXTGmqz3ylmPoU7Tu4TIZURP/95dqi3BHf6QvnUPTKGAl4uafN0PLzeEkjspNN5/C
vni04/K/QKDpgxa85gtsasDqyIKmwUwKZM9db8gdA4mIUc8FLdgw9dfgKKI4tgB5EpPMO/Tj4lis
tqjm7rIoMX1dCl02nm+cc00Ed2SnpCSRajJwqkmgz9Uw6BQK5BquKLHcV+uKhZLq96f6F7NxXbnC
VSmpjLjMAEWoUhzZfYGWzNZOcaJaQoYR9IXGrPsoNr30J2p3o8wNrqGikw9KYNxK2WvLCY9Mm7xZ
ANoDsp+v7SBkr8eLvaW46it+Y7rYG5klsRcSUw2nGHzcpwmn6qcJp532CjFhZ8hmxQdCEJZIwILp
uVzRdxU2t90fe9mLoXkrhCopSuvSplsAbKZ6yaOhsSOu4PuU5VUVh/u6OF/PfBHMdXgwxU8FGb0y
hUR83gXciXE6dREXeQKuXfCaGYRt3sEnSdXhFFTMqzCvmb7EX97OWDNl2ogFkF1eh8vEFp0cO/9x
ayCzUdCED5U4SZwamqb/MDo9zUz0PLFfyfocYTFS3vlN2VJ3g9+6zxksTm1dsSso6oHVH8ZJP6wd
KIr9m8QKTd0FXZnWiH8hJg6E73Ssrjj1b7gwI40w3m+jM0O4LqBgHZctjoM+4eYsfe85yhVIUyKV
Urgl0O4NuR1uZsW1VMGVtyngNkI31gbHIWv572fxN4ikoANmSxhGNAG8/qCWyXdQfJUNELlRqqQa
kAwhWwDVJZ+k50DJZTz8jARz55BNIjVR8ErTF/GuvisBZVjiueUM3GW1QUQeP/jr86MB0LIYNccP
7DHwyT47vp2fhU7IuvD8FiP6/DegR7eAvpv3T+B+xcT/I0uB2x8fDgPJw1/b7F5HfvZCIbNb5SVH
Tw7kBYyOuTrwFrANCDbsV1429WaRXUdBnqS4UbNEGIFXNSPuHpR13Ge402Mxb5MyuIoWP6pRx+Eg
Pj+pw3+oMLd+I+j8zxN+qdK0FuoI6nIHh8NDD61SHNGXSOeWuJ2wEGqziBE6o/rm7lnw/bQdqxSR
YV5Byzql8lSKdW32uiMMYz5nKDMtqxStIVSJkUCxjUlJ0mnGjcnXo5P7leZKY58LPiS94oXhcC1O
kzKxrKVJznqpGM6Eln8v0BX2ilCKY/b4oLhLU3B0u+qFUU2olYnVfQhZM3E1Tp5gS54P2pdf1v7c
KMuRwNntpy+X5hZYMgazx7Dov2KLO0FXoYNaiIj/o15wKmxexJw2MwilFA9cGzvh4CMHx38XNzKc
wbmBHeWpHQ2ARcOylDwPaiSrZ5E5d47fg7raWfP4ysjybfrEWn85I6dCXk6w0qhPvAXOiW4AZ3bh
xgXiJsP7o766J5nn7rYPh42eWEfuBRnR8dh4lgEAHrSM0gB69R5KiLHVQ5/R4XG1QSCw4SsV5Wuo
ths/6EB8J3AY3AfdjIkHCCeVbt5x8c4K68sXKhTR+ifR5K+G5ToxIAY+OhoJ54flErjCOsmF/Wiu
rfX2Wa8sXm4npR8kPiC5at4zYcE4qRzc0xiEcXBo9v8uBV1Vifu6gh4z5HlYIFA5dGnrDkzIlSIK
dYpVB9FND7PXET8E0tDhT3Flaubox2Hq5oXdATN8WCNhrjM4V/hELCobdz326sZQhR5GUkDcApny
8Tu4F2YAlvhn2A8Ni4Rj3USuxSiyNiEg1PAK3+1XmtcJjKSIl4wJRNu3+Jr2xP+LlOpkl124rb6J
Je/Gg5bnxJndk1c/DuCX3w7v8cZrwLv1uAZ/6bzHmHGswjZVzzR1xNmjDtRzChlCNkuAEz2kRbLx
TGi4H0rYWZ6AR8ZksqJiY4ufxrQg6Ldr8WBUJmMvtPmytfptUDr2j2sHyxEQFfzzya/rhjL11VKL
N7QNG5cVC5N31XO+mpdD6mn8gvddDzOl/qRc6SuOJsMjfPTbzBexpAWrLA9YSaGy/2R7d9hDZvWH
f5qEB1TRWgjyyKuu3LEVeIMTJgnHmeCOujSjgPByFLXLpFVmjFDrB5Aq8cu3WtWI/NfA7Qem5gy2
xsEwm5qpaMi/nT+K4rQPJ1N4gMikPiIoIGI1I9NSxhJrh3PeUJNOh4qrXWU1Wu/XMKwZnPCe9pak
HvHKNuIrD/jHS7WIas9/1iLRBIonDsenldC2bBC28pf5z3WzOe0WPpYYaGQ827RaH73ls9i955f7
qkA82W14/tV1nEVK5kYtL2JaPDbUU6Mfq7liEafhvOXdTnHAKAykh9k7HNAniy5DUH0nnOe3lVjG
yr29Ha3farSkRstToaPVDiM+kHJ8N+TCwK72uI7LbeS2+2LQRlVmYo4X8PY/ASciygc1olGkqFh/
qMNFN6cO7zZhDXiCSeSPwyvjeZXiiGBoH4a2w8IBU2AX7tG5MDMkudV+spTesytgJcAiQs6CpfwF
XsaGajW8R6h291d3smw/AY5JVSjZsYTSvsjofb2Zxm5nd5iL3iWJXoeWWi+3mZQGkXW2BMHF2CVS
71igJE+ptLEY45GJad81yapgU4axkimT3BMSoPqNfhxO5OV3Ta3odZgdYhdqnP+teV2RG/M2Hd/H
E288O8tfTHu90FcsNy/SgvOzLmoPcd0/jHLd56BDI4zowvJ69W1PZyNi2AgFDDHSY64wVDAD0Cnc
6nomSA019TnER/cjplfR/my3/bQV5gcWPTh84/J5wculwphZJOuhElTGmOEhV1jeyaq1Fd1hzTTs
lDb6D1sOMQmeA+lhr8nVt4CThr6LEBDzR0DwrW6HQCfElBCaWqCbnWiKiR4gJSIGEzIn1YHKLcCu
LfEe57KAA1/tUdDDJawHF9BsHlIPOdLTLTORxyTMSOspPtX9NVSGGUWnVvU8FmTNgyVplcWAXUIT
ee9Yg1GI27KLGOkDIezcY4sXmfonRF7zo82INxyaGwCGcRsv8J0VnEuBiejsOBoyo/8OrBH107B+
4mAc3+SyCipuEv1GGPGUbQSbUFhd8bAFZSgTVO223XsnTnv5ewREPpjR9QrBsdWdEKtHRSxfwqbM
mtPlrN3vUor4eQP8Db4NpsWWkzKRD0rVDSpXhpK9d7HGXIHpk4SXGSM9nTh2+e8N/SFKI9vr5mx8
NwwnSy4d0+wgkNtmxRUXUa3IiPFHU/+hE3CDn/4ntwb2GlKBRD6Ae6Y1ehUydDMTz38WN6cs7mwv
juVogt75j5Nk8CmgaQMwbkVFALve36moW/zZokz4L7mitltlw0/FYgtIAe3hqBryx2rQvWDf0C2W
Oh4lru29HTO/+aYwUubowRlHDa0/8At1XdjjdkOuy8rdPtGqpI0CZAJ7/DqNlAPa0gSfKT5Au7kP
YjYpg+Od05YDKTRHtEL8KTagsyy1mcf6P7W+75CEdG4k99e3J2UIXN59F75xz37cnfNt2zwWo8zU
slA09I2lTSE/zMRFXLwpUL2OZTCm8sTOfJaF59d767021lvzPdEnJkGrV2e0U4rQht4rm6Nx7NfE
Ki7tT5Rhe7FyvdRAxRhjmY1/2771QDsWk5mnuOrc4cZz63aJ/cxz1d4UJNa7TDqO2Zinpr3SbAyb
6HYsI3502PxmvK5mWOxRhmbtA5dcuDOFHSCvJkJn1Fim185yR3CbSqJ9mnavtlCY+W+hHZSUVg8P
syLhpJ0i/j2nTpJ39m3cYrFYGqRiBRf3ZDHOn3VFxfWqXpo8WCpeh2cm2yAL6Q6FBMulgN5Z9gAt
oEvw9gP+CTbAiLK4q84JfvUWssnxx49+USxDBjb0IlqWNFGpzv/JQE1jhgELytU0IsPHKFXXug8G
TXYg8h/HyNAKbpnhDyWmCJTS3Z5AfwHCFT2u0sAhLQaeDVFw2DU+IHWOcnkSfnbHElFir4Hfu7rd
EwOcYOgMs5rDiaiTrZwFkK3CKX/1kyMs3S9IgPKgrsXz4uIHvTMzZ3hQYXTC5Y4H9cvlN2Ax/ZRC
0W85mvpe26738kQ52yzmvf7eqJlgl1cNSNii+RWbbZPbk3VhTri/nlMmnwYMbD5gjWBY33A5gqfO
sBDn+F2O6Q6rk4M5WBHKAFleJJdf5IKSkd59TUsiDZvr1UFZCv9Ppxt9L6ZMPy9644PmqeX5TVzT
YeOGylwSDlWtAImiUHOWL3hxFR3XPBou7REWQHnXkRURf+MCBbhOauPVdHfwNkry3/ByP5JBD3RO
0BbSaWAc1Duqhmfy6me5oniY/6iQg/rrtyJ3ZG3U3qLgExk7tn+qxHRVV7sb84TCUojRsjdo+DSN
gk0uEfGVS320FuP78CH98RhDObVqWkjsjb8HxVbFShRf0wHoXjGIYPvSnKrT9VhN+VQkKCmUF7vP
48eq2mtrbmbOlfdkVMSDgUjuMHKhpN7/X3gKEQRaB8ai+luUtEXTKgF6vvt82XMOTswnQmanMgha
0ENrZ28dHSwgE0Snob5mYlafk1QsBazL9KuWopmgb4WsXVR9HxAkysmOa6QShVfpMXgF/lurt2eK
7zG9GMPp+451cr6BwWxmWtN9F30ZuNN26EV6onk+WCuwniVYsXJu5GJl2eATWA7gT6yNcwlnAW3V
N6qJ5Ce802YxQyYHGqr/Dv9TRswto7rNGkIkpVTE1D4mO7zyr4Vby1s/0806/bme07JVbOUotqbC
SVbJ0/W9m8tcKHd8jguDPJ3Wo2Irur819WuhbS9i1LjzNjsckztEWJKcRuCslVYfcrM8VIH/r43M
WxzbhyP+bCshRy7wEImhKIWowgsqM2NUPjzM5GY9NkDtf36bZmYZjvqyA4iXuAy+I5eQKVykV3GV
nd8rbTqJMumcSCIoB8T4EiRkEdX5b9xSrpBVOHyMv+LYnk59mP+7w8WSeDfjkIGuUPpg115vexWa
3mP3L8c/qh/AAL+/IT48uiO8fyheRJ2IXCSQwe1KgTibe6qeCPLnPWg9OutX7ZOENh3f3C9HOPwc
G/Vdf546gc0Ao4Xg9HiXlbk68HCRbcV8SrazEXi3nomQsiTxjv3ZDOQT3yZREypy3t2lJp39xG5e
x9kMEc5NSczN3Sy11zER1sNG4HxEdMYATQaYUaVp7gctY7aRUFeQLWoWulNSVvS7+GZOeHMkHw5/
yRlZwGc+cbBTXZpE+k88139MNA8KTFjmInQ/pSK4gRsUKnOSChFGfMyVoxV3Z3603dBO+eTDGCIg
sqkfNZAlKZy4ewZ3IDFw1R0HQfctegwFKqK5k+b7qfP8TbB9CPlk2XYNoaQ4PV6fKlUOZY6lDZYZ
DaNuEsxmvI792YipnSqZ+NyjfOyyCpH5DXj09Ol1XKNESmxOzpsXSaHKJxV6Dz50wZl78nfMA4WV
uJnsePvE1g/OGZaDFZX7pPEFBcHzHoQ7wa/lPUlxhTuDYaCkytVl19ZJb74X4yCD5SCY7eLuOZ5J
f0zj7uwPjnLMu402QSr7htXY78j0+MhoC7zi5vUVBeqeXvw7vmsp0zxaghJ+DGJEFei2+ROSKqSy
yWvn3lU+b2GvYmpnTWY6XB2MAHuAriIgJ4ruPQM7vf9Xvmc/GolxsRVr/t6UH4tl+67q5X+Qsr5e
eLBG4eWagKTrZYhLeeIhbsYG1ZuiOGJYVIub4e+StYBVEGtCfLzB/fJAsRESKF982kcbeg0M83t8
3UYhH3o3OE2vQX9ez+NRvo5IQF+wivGT0SK55QeQd/fRktmwSBHxIiB1hQiWy+GPj7hwHJs/SROW
8Ul042DLYuUKLkfgKNnWp6A2QkPGvgTaZI5mD4sU6okw8hErv3KCMrtT/DTepa0vSCzaZkfz1D0n
0/6wdQ0UNam4BKxH2AC8FPyVcbOdzlZNiNLUGjDMMIqoqDAJqK0y4gykOMgBn80S97VestIWSCsn
AFFReSu4bCLu3XlH40qljY6wbCw82dEgX8zInQ285Xyr9H9BnpfC0yYVkuNTu5a8qFNVEpc2FW5N
1xHep8yYN3nWEpc2EKdOzDiKYpOzXlsmrqDY4lgGiQHKvHzYSMzlBUgQzrr/eaKeeBcg7lTkXIS0
uE9xM1Dnxrjz4/NooqxChQyRsqNGIxGnTDEZkkNesW5drt32z6ILExYiTPVzNAMKMkWPxLrz5OZO
/RDWzzMteLKyzGbRrbL0UTJqJ7KzUIFO287TnxLWQhnmk50OZ1mk/ZPWebYjtORDeQ/ksyoAcsT9
FOeAx0Wg/WUpMjUC5rlx+9nQYQ2rVVQ3tPe9GnH/AGm/SFUDvpWQ8MYFua67HgTCbEzWJM9796Yg
xff1U8MwYyGKMajYwTqJCx0LvDlAZtH/s4Bjab0Gb/aRN1kF4mE3tO24yRC0DtRyGX9DV7sx9T5b
5EghNagRvM0iftiYTaeJDEKZ95sx4pV1/ITAzm1qeoZad1ybAiiGeqmAzgDuciavuVP7TtuMYiGj
DqxdbI1ay1UVo/e4DfY1Y4+uu/EtFj9DLXKD1jeEtkYPgzgKIW66JJarx/6BLgZX6ES5CkvhU7ja
B3FWagRY5+/iYjRPL/R47vQq/g33VIn6pTp78y6Ez/uUv+LDfGe1J6TuSdZuvhNgyeU15VnRKIym
Lhnm3qtqfv/angAozu26sbPXYzWb38h4dvZGwUZVD/a23013aRTClLJy+QDiRaxeGgF9bnXh8jfg
RnCAYeW0qRvv2DgVRWKFjUGkJQqRfO+wMd+s+iY38Us+wcTD4qWcdW+SgY+7gvA9R60FA9g2Z1MF
c0XSHj2NKu5vr9ztETZjqGJ46nkpduHBoPL95u7CaHDfeASF6yoWxgLbDswJkfLuPAl96TfeSMFL
8VG+f0VSV1EN/CL92AQqm0n6KczWCu/SLY/8PmY5sOTJMVz0dvRyV+gZBbRSPtixs6eklHCOMSzz
pekeY9VydYZEqQ11cmKULGF5/zNgA51lHjU6rRWOoxTRtveEyLiPz9F9zOfSJElhHH6b1R+MNkX4
WnLs82rY/3I/rY1nTNvTZcvmqGURL1GdHLE/c2WwSmWysp6hoitzNoi9stuE+6IXnuDahIvI/Paj
AjxhUbZ5TxlFZ6RTbaAaE8wn7jrp8wlBb9KVfw8SliiEYExYhdbC7X3zIr4+pR7ZDfxA/sbWx2qg
IjSSJkCcjuhnvzdLHBaQJrN1HmNUHYSQUBL6eolvzAzISiAdRNbDdJEtrYD5xUysTi1SMvSylURB
gWywb9XtPlZMnqMPDgNLpS8iL5zbB/mHbQ8HnYPXgHd2d8ecCLMKVuyR3wrU+sheD6NsAM9E1uL+
w86Z2P1C/UZygh3aAzBFK9/UHMAzM5K1LXxk+Gebn4AyFohrdVamFp/cljywjlrpVqFC+e864pGs
fuC1ghoEq7pMFhUOiiLDLI7tmw91bX51OD9hnarCl2zJmpjwLQ4dIKkexZFNTilP7hI7dw3HxvpS
CmVns1GH6E+t
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
FF92Y2BScS1tYCbOJ6nl/yrS9tO5nLdkcinIUmduQUlX/rEFHoa3Ivyk0aB+kXloe21LQE4kGkQ6
Q9+cOvbtZsLXojH8eCz5LSxZZmj1OY0HgImQvBdW/AXKvPSh/8qp2AkQS6z06aDmakr4JM27sgw4
e8FcV4tuRcqkGs7bb5nTeggXj+gCM8w1pZjupaF2huj2/7utBwg2caonPL9QnFqNhJnw1y8cEijm
U2tA1t1pCHmc/cfMmTL1KVw5knK/j+GUCQdryhHqwEoaWgcU/WsJ66DlhJyiBG8LqQzPrvznCBbb
LaJ3ZRAbBz91jljSVrMpulWLCnotPmY5QRPBNQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
cqAgpvQThUsKP1YQSQ4a4I/shkrWufEhsDBDReUcDIwQgy0J3zK8Xf8BMFoFrewCsS2KNDRzQ+ER
jCDGccgdbKH/8jqChdozG61idZWa0ns7506SogoQlXjlqxzJaYEQMyNxDX7Ycmqi2PkN9cXJyFzV
5txS0QofbL3mzPtdA044rsuP1fkQj0yHft0ysK4zktjTKWnJPMDoc1p9qdrOCvbt1ZBLB18dsflT
y4tm2j7ie4QPZbNefa8AuI4j7gxnCkSCkqJB+CSn4ks4ndlDn/a3c79q59d4UozEclqodJLD4obY
Qe0wLjtJvGaBIVSj8HG9RNO8kRI3GFa3bHt0Iw==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=38016)
`pragma protect data_block
GMWtVErQpQVB3QwSqSu3WLxWBruia83TiqFim1P5yolu2OZ1WaMDiEaix1fNQpqppRVnl3TkKEa9
vcJHFKzyfXJqgO3ZH3X9Vd5QCdyVD9cyel4/qof28uhn5vJUlmrKomzrreR/9G9xiN7OSLcynfnd
YpQHYBrgKHNXyDABRyEMAHIVwA6rFCQXgw10Vqiuh9yY3xYnPkhfaG1ADOOQhPlUAFVHCPvwxUN/
9q/zrB7c34w49qMG9AX8pkcFKSI2Bf80mktBW0GbKwCaOuuroKqhBP1i0QEosE2oOuZs4uznKrQV
pUYsw2IBm1++2cUcg4e6k3n6xJMjPgSMAEhoW9yEngeVWQcZsBBAaN/rOqc9CFVqP+46tp94pmQZ
b1w9JLEnkaUu+UlNbuWFZCCTKgXcpQa/25PbW935TuI+us+1mfkAB37jCGBvh76OUHx0vR44T4+q
PoDdHQXqDp0HMStpuaanvbG6WyhcfOMiK8ICrMeskteftUnBjUhJWVs66JJojnT2lqKnSJlasg0Q
fp4PURMTXM5l9wXi6563FDs24Nwg1dbsv8kCSS4S1mDQM9EjJZyrOjdyMyNybw/LgECF9AYZRJ2A
L1PnAzXEjVxjAlPH5awpfmD7jTtNfeE5qXMEk6OWSrl3ErXoSWjBY1L+llf40S3AVes5uZH7scSi
X39jIqMklw0PSTwvENkxiQ4Qv+ZrGq5/v0hrXNA9ASetnnsn7C5nJaRkT8lAgYtMzd3c3zucxfM0
xGMENBQa6wExqHYN6DNcZPnpOnlNaCTtGOPZ3wSBpNe2WvB4McoBIwDr4Y8GYb6GO47od8veeDUW
wB5iyLW/DDKLe3h/9HVLsR0V+JWD7hvmTjLPtm/89V6j3UZ8qbUGuG0VOAuk7XvYjMSJ3Yc+4Hhv
rZLhbvbeeGj1d7sR4CENVMiSh3cxBz4Lh1fBGyX6L6o2vEgE66EM/cT9Wko+KdxiynKUMmokuG47
BRrfT01g+Mt8oZFQ6Cazixd5jRV/0LJn1OYEw5bKZVJdDAr1+F2iDl8DIrOgN4l2cMoPtBK2ZqEo
ASLWE7WY5QpD5AA6OpmXI/zxVfO68/Brl72ObyIeWiAQmWGGv66ERTZkQa8RJl64Eog2WZGHVfWx
0axfdir47kWsDAL3uIqPOz1NP8axA1EKaxB0NR9CcPxfjHAjEZ1T0fmk28vphw4h9s10ObFZMCWY
sR41z/C6bDli/F7J9NE2IEtfN5ikTtMNGTn8uvpNffLCpOHmGnO1u7/CCbGCpb3UMStZPTs50czw
J9hntiN4KyQje+dRfTuclk/xKESgQyWiE1+EHbITZ8iU6Yp4NBVtJpCt5Fc2fwC7jE85+Ptp3zyU
ALyxHe4EHpGEtzwbHtbpg3W2UWEp4zzMPFOE0h6nC3i9HLh2nMu9J5KwbfM4LGf5mP0ovfA9zUMg
if6s0TvMhCbAkGqK7/FOKwZGjelCNmxCoBKw/5K1trxRlF6fCqE8NiEzg7CvdyHgOwb9dSYQT/WG
CTmj7zg1TCsgCe+kzhTxJyk/cXHuhD+RETDrVLigD1Qx4D11NiC/ve3n0wpQ0gRMqPF5YYObquCC
deMFPan5anqKuQbw/S5lkC5MoZCvZ8BCVa0nVW9bVcx1KWVIFzhTcZdxpZT1A0wPqnMw+1x72N+5
Xb2sj/ORqo39PHA8yN7RQFcR/L7d5IN13Bk7K3hnCS4yobHpCQUZAfo7V3AWJfVAnL2VKy6wkxQT
gG/00zShKC8ElYtA63aEmnBgQA6deIsBH6IJNvVOwE4fVcqj9wW76S1/Hjbm+IgO5kt+NtsMvOMR
cno0wbWQVBT/ZoXhGiCr6cLsro6L884m6/2KLBeRW2f73OUNtpEvF8a0dNMNXAy4llOJmkRXeVrQ
sjdl1XkhvyEpUFe4Mo9qSdPsKI5yxuKjyq9e1SV0IgvNkseOz8AFg8PPVaq5a1lQOfmAiiiltrp6
pX02cbSJf6V7ldoMd+JPL1J/A4oae1stPU1dJAlTV0berEZlxkcq/8HmrCqsfJDHNfuZbNdg20P+
5xhGe91/iIsjr/dqmDUNSrPMJrj1Bj3oKP9gxdQToLtwmldxiigSi8QlN7JRCpt4X1Yb0jYF/HCC
L1YZ8MWrODKUw5HCgFebuAQ1Ho1NofQoFveRJRNnJR06hmMAjkZefIHmMZYCkznpfS9gg5MQZHDr
N496VD98oIFvbqrUPwaU3u6Hr23S9XjtlH6zccZHYVb+008yyEzMSJzWSDV2mxqEBT2WfKNTxm5k
2wDSNHxgxSiGYykape8u6cg8OCdd1GChrLoIfHtD/qn+nFP0fur/oFCFW/wzGXxuTEvaUslDJjxv
N87M6JTDmhd4LC4m8pbVrZllvjZqLVv0fKKolMdw48I1AXuExK/i/IfSU4+QjPmU0BA0UBDVRgM5
WhQp9RwEnnHCNr0oJ+LjddsRiw4E2/xBRD0oSac13fSb07f7z5+WSoDfVLKg2bATZ8d9yQkCw8o5
ueGba4Y8YuRPv94hEOl4eMgXeKjq8fKpUzqVYRJa7Lfx6nZ4JJxiWzZz1g2gtIlpbta4iyewQecD
oaQqF9IntL9BNSG2a3LzMIfLeMwcrbglSmZi9nqmxXDy43qgH8G9VZeaQ1eLXXU72fTuN+ZMXdxx
yNIOUEGVWN70dl03hNFUk1VA1E/bj8hx19/5mNrAb5DO1gHrV0+/morY/e6v0yh6GsBQNPMjVTfX
fTM/m5h1aCZ3FFgI9Ae+B4PkOGT4kCfb9p5QF6E12xIDIAglYjj4Q1+hxuvfh7ybK+4ra50y6tzu
mL60PJQ48bEiSgkaGoraGCkL62wz2Bs5m/BNwERzO5eW02dVINqYCQ9tXKTSKXVQ4iuvgapfmFfr
Z8ZP/tF8ouaBflrH+rlcZNk+X9GKUzGYMhkoSahd2khfPvOGw0uLE1dbyhUMmnpEVao6i6Xi7c3y
Q+st4pd97U29ae87iXfQweevAebkQlInu+npuPeQx5gAjfcjdu+AJBDnJKlzrH38zYGQVVPjShxA
VJ/+ADRFUJf/bxdGq6hl/LPYTBRBDbbQEft7zwaAnt4bvswU+GE9C3Ut979+vKNvqSewHi6WCcby
Wowpbl3GIz1kjgsRbOIntv6xvdLOvKqoriA6Khp9dxdyU9IaIcS4H5Wul6LiaPqeDNkyI7WhvQ4e
nZ2TmJvpfG5ZIRACSlhox6tmPl7DrUf29xeaqsn//+nZRZNRT/r2bhCqQSrwEw7vThFHF7xxDb92
HL4U52E9fVcxNQ+YDHikgLMnNXJB6HywTn7Z9h38Zvgf4vSlhrJOORlpe4raSbWCcK2aV0XTmJB4
kX5UHcu2iDQ3fPq7/b5PMmq/UalK/nXi7v5vwQGv8JBfjS1T6sBfG0p52DY4lNFZs1YjwLYOUDji
G9LpRJz5pY6S4kyrV7MafHJgTjs3gNFdw3o52uzV1aZoWXNUnimQrrRmi06Qao7h3SlVscR36tvW
Eet+DGveNy0rqSRrZQiJ5i7liH61I4Xe96YSU11VmGGW9Rl6e8MXa2cZS4qvFPoSYVrPtdZbtKaR
Fa7StwZVJKaZj+D12n+lBp75+h/hunHcyBeZQzpmmDVMjjlnaFzZ3E6+PUsHrNqFkMw0qdjQcCew
Mr+DSYXQGj1Jnmcu8hX9KDSSiEaAPA24om/rvMZsHw11g+dW2JHhtIqwSyGpupDz4hcbJdnuWxcZ
Y3TYcF037ehWWy2cky/5rJ8NBVfgsHPag1GanjZK3c0tM7fm4WpKqDkKNLGFTaYQssAvztl6eO13
AnA6plQXvIXpc/oRwaf63Q4c8GltU5PqBViCAHhFd1Xh/oSldZ4DljdAZpeys+5gCgWN+ctoKNyo
vVJ/SCjYXnGQhhzCZ+OZuQg0tORh2N5LP3vzbtuHmA57oeGzKnXRN26tFBnVqQbnwydQ8DRGi/PX
oSENjkV52hRG6gxxiz+kjIzgM9v5XuzHpnNO3VmIT4nq4yxeGvXluxUjmGuTXjPV0Cbx/L9ZrCvE
4B22rFeGbO8mSIuaZ9Ct1S4EVSJM9llyKyZzEdKPuaJ1IScc69/srMaj7pPGYt15h1BCHEbmq8NL
nBuu2W9C4kbqr1qZ6/y6Fj0zf69CcztI5re5194EtqqNou5iAUyEWp92Uc0aqRPG6ileW8GqGQQH
AHZ7TGsHjJfwMPsU46daze/oyNItz7KgwM3fBcaehdM9ZnzlIRljeJZ+nHXV6tqhy26Zsy3NAiEM
FUD0nELtBqhuV2UOfkVO9O/qpZZftqfyCihtr1xTKFnJs0RQhXXV0SVzgjAw6PinhASN13WikEiZ
slWcExNXG4ANWSRinso1bWmskR8g1+CzPJgd7dIZRe1UkZkkSZhL+y0bv6UWn0G20a9jN7iFZJ1m
gEDdPF4opU2Zawt+ogyxLqc4viPVrNDC81ldw+V7c29cvIu9MK7KJZTbq3mYdbyKFyoAlBqUfBPE
sV5w9C+wN6VLV18tqZPK7C33xyuKb82l29j6xEpGYnS6ssMsBWUVk6jaTXosCRxyDAzMfHm8nyBw
LUq1+gFGXjU4Swr0UYM1uThedMAeZ2eOqtNYvsAMNU5x9PUoJuwLhA+NGiTnaVeL824029HU1yDC
/piCZWc5J+8Hh3qle2LpfpxLIcUpiXJjzb/WX7dJ79nmx6ikA8k9ndSuhd4cN/uSC6mc0TDugUqL
htJnCn6H8oTkZXH4TTtpWLw5LJnYGEgwMqtoPC/n/7llBwQC+RevE7RmUDwnLPqIzeZbdAYcYHl/
uS/dWUTGZmvs+hxJoVl619u6EdX4WL8jxR8SwBeka0gkYC9+Zk05GMDMOvk9LAzODcWWe2lC84AT
KOO02mQWfVqKF66mRjd89OdJx8RN73C2MxowZkzTWP6xrBN7dHm6hFcfW3dnnz6SK/uFZIy5bj/G
Of6Vnt7Hoi0GdiQ0lWxRHLZROUv4AsAFSZZlUZfFlXZ9xkA5tT64E8wxNln/XfvWBHomOSmuz6MG
ZNvN2h33VsBWa/R2KMGsNBLF6qAMnalrmChZId3djg2CO1qx4wK+FYlay2Ud8xkZfJGNarwACWRC
/D3L9r1tipsr2oqbJ5T9jXg69XqelS7p2Qh4VHo5Oqt4dEz7eSb5eCZ87gPGUqB/bRNcd84KZ/O3
rZRfT7GV7zJ+DXYk3J2MUqI43gE//wBMFlSFKQQ5YUIaomSC3OROFVIbwFAm1XgwxkPR/QInsNg1
8WR5NgFQ6Qy535xlgLvVwPjwCXOYjokW8Cj6CZY88BwQCUyHBpSslox5/rsQYpndbumwUdHgsyWB
jH2ZWci74h4w2xbr08DT8V/sSSvywUaA8dIqjG/SZGf222r6Yga4sk+GsUDkIwxdhLVy2Lq7hIJw
DWy5LIwNM6Mcx3c4YP+aasQFaxOqokmtGzuWmR88Fs5pXN8Dc9CmRnrRFoQE2sgFeKmLz24K9BqH
q4JdG3BouT/p8Ty2NnePF7x4t45DMOCObbmOtKu9YAVrHIiR4YJbJekzNiWMgJJPgW+UW2SACa72
jK0q8SBEyQSm6tUoZnLB9UmIJ8JFTml4aI0sYn4yjsAm31jfk9Wp0aeUke3Sz1qBrX9hwfbPSF1G
Jj9jEyZUXHDUHroV2pZpZHTXGwOOiGsYBCmspEz0k52D3eOjyf1Wse3JfyRCgUc1Df0AQ1nC5/w4
BCsE4nFguehLkVdbTqKRLWGAkhqj1uMH1Zx+8bJGmhy88I7Gl5hHVaMLf9VSes0ztU0jGcfeAEJp
AHLw65tGszrq4IqMh4haUY37p+/HDPeQpdHiKgXF4KJPamvMq5krvXIhpMI7w0ejknLIJOQOIgCi
CJUvg23gtH7BCbhNsq1BnCOIAgcXT/BjypoqgfVSOCMyJkvcDGJRbt3YskICzpuMDZ9EPenVj5AC
rKfz84kDrTqA0NqSyI6c2vH5D88wO/GrIgyW6cV7owVbe2zU/qPasdGH5r8mvL2VIkp9JPCsV0FG
JahBfScHNe32Zv9/17eWGO/Zv1ANWXFeFNaGJCAVuMZJ58zqaR4/xS+6b8++70YUx7UUtCaDhYDs
UD7imaJsgsfl+JW2zfWcJzqwRcwm9nlK2XCDQgQYG/dRdWWWO7E1YFJplJ23m3dcyOxtEnsfG68q
vLLfEswk+xgEMUvpwNMtm3KGUURUycQKxK8adKmD2mxu4M37KPIIU0IhOUVT1Oblcuu8aBlpls1n
oa6861DsoMaQ0xhFcaty8sAuAvsMcUcHLyVXRGAXtAjvsYQ3oPR4k0RSGC/932jJ8w9lme/M25UN
6fmjD6jS7IUAbA1+nPXaRtF3/R5EZxH8rM5LzSNMxwY5JH/On4AUV0ZxuGjXap9QjBXE8IvgYuVA
vD54sCA/lGzMNYTHWb78xDfmd9bd80WlvgRVvyinhoRA/w+c3BLf0tdiRI1YGOFzfug6Hxp4qcp1
blcrlrrakR8ZOEidU+oBUI9Z2EMgFe3a8yQA43rNAXytFJNVcSFT7R5XJ76SadU9dyryps2+tC/7
W9xZb5ATscBBIu+8q4ZbzGQYhBwtABtQxTt9/wKZjhsG3b+lB/wXSHQu9GWlgbHkDqdjEg6GwUPd
yqFXHmGFF+Jivx9aZ5/j57RzBXVnb18y+qUJp6Sjgolqjr5rNqHAec9eSBckqXpQQAsjAqkFUqG1
ibi0a3Ka3OBNz8CK6UZNSUQPFJjhQkAsaJ0OytLaKICmjo/P3UwAPqrMY7vV7AzUWS2sJ5TC6zBk
ioxiT/H0J4zWkl8j9XCbZ3mqdqT8VZx92iV+IgcfR/OTaZTJvXDo6DAum+UPmBxI1i9EcX63QGyY
kYNGscqkD5EExp+2qkWvsa5G9vBi7ZJQ0QM/8xz9k6nr7F6RTOWwdJFbGCOq2C+VxOxY90IwdW8h
HGV/XjGtINOvn5XE9f4TYESeLxitCv+tc2gRqrZuTJjFeGmyhvzbCJnqCmOm3DNLzRiL9Fy/X1tg
ivDnt85GX8JxBWHNmimkwB3/PihTRaRiKyVvzKGkx53LiihxoUhz7ZLFeNcW+jDKWvB5c5NviENX
/JqxhK4hU3sA2DhMCSYXlCKQ5i+lbA6UdC7V1c6OXpCbAWQj/bwuVE1JYMN7Hm1+oIQrHM6S5+M4
ZiXXsXcII7QQ7/hrzNY509hc005k3L6Ib/hAoUwWQ57jmgQz2rZl25S0f47qmhzvrJY5gmYCW1pH
WkZpI38/UYDZZIEvDAANyi4lpm59v0uPIwM29DkGcZ4/y95z2LTdxqvzr5eLUePMrQ0Ci3waKLlG
3gVUN22hMJiHSiDQA3YULMug6UrCnvfLKnlK4+b2Qz6NkUIilyjKHzWzDtj0DEaEzMmsNBFFaREd
VcQYaed2jIcYwd22GQaVXKRjY8ZmRt77xBjwXlI0av3ASjoNac5HScjz5Id544jnPqXfp2RsYTaf
c4g1pOFPmI8VNrtofpz2IUeM6ovIXVCABEANsSCbu9Sry4V1mTCA2CvHpYF0D5CMTlvablXR26br
x9XnNfH7TIkJ5oeEZlhrhf9DhTWtFkFljiY1wMk6XVuYnn1/6Q9164++46tclScvDiFqJ2RlmygV
83W5seCQO+8tEZqrnB/+T/R4zMeau83Ah+lQGBqofF6T6t9t68zG/MFADVcWa+X7uCnxpuD4me3S
ancuCXudpEZ64z7Ykl9sCKQyg27Fjj3+CmJVd2S4KUjhJUGGVKuCe2fzRiEZKCKT4gnGAJDOt0Sn
DzkxmjU1CIOKJ/vTb/jCasbo5OWBdL9vTSY3xsQ0TH91Q15jbPeEFOxUh7797mYUn2IZhqmldvSI
RCtqkHbZD/l+nBHKF2f5c2bns/wB9HzUgrfPGXdA5W47uwh99ANQTXlHSqYuY1DZcrGBVcAPjn7h
JCD8J/1ZRi7FJZuvvLjpdyZYc6Y7V6n6Q+eb6z83KLxmFhfqQLTbZuINMftRNSKVts4EUiHi72Or
0QEqihuqTaoKwHaLgxet4f5uLVGem7taE4ogaSXpR0ipJdwmE+fBuFIr7/Im9SzVX5sgd6h9EgzZ
kMBGlTj9OtqHR5BbM3PFEAgjJWLX69J1QPZDztyWLlNNO2VvwYpPLvMjNO4quEcIHtk2iqQQ3nyV
dBLO1w16Tu+uA4ghq9U0dYbBJWvMgfLpfTMuUrzEofDZb7KVFHEweYRNYLAcqQxDwdWB16M7svlf
/o40C/xzlziKW1HEtsJX3f0gwvtKYF0vOuyty8A+MkyLPUbdGlrg5TlHbMf7/chZkF0nB1RGkmsV
uCBxxgx9QFoWON5+H8KHXE4CWEvyzP/oas3Qcicq7Pypbqk89BO4VOvK2GcS7WyIe3mFl/xSGiqK
ZoiukB1fr5tNcw3xLJwTxyb3rbUoDZbEZe7+BjMxACNI0/IMuzqGibEAPMZB3FMZdqn9aPt7s3vd
fA8pGQwYTGdtPwU2MsvHyT58IaBWVBhinL43BeWeWiiAVW8Jbz1gtq13zXlacKVfZF3y9jjLbsqw
MtB0w9faBLLLTLRKWY7WjqlYMaMyx+aBusLrK7+Rsx1KtQelr/AkVV5q2uRoIIjknuxN7vMg8nPW
1yf4aDfU21HSCQ6dL4xm/wHzntv96EejFdDEfobcpaT/xmU42Z/SfMtui/R08GG7FtomH4n9I2sh
LuyrIV1feaJ6iRtwbgtX5WRHonLe33gCSKQ9i/x5peJOiJSXW0ukAUDTreo+ZzZGUQAPlPVlvN8z
1tcRx/tuVkb5TAQIaSYtMJnF/cgE24CstwLM2xXlUJ+os5ieuJc18G3YCoevya8IDP0fQo9lKnfl
qQ2x4gBT5WwJ5f06mXG3f1PDmNpP6H7Kqs0jDVGDkq1u+9JWXLf5XG6UTk2ipyHE6bMb44D32JML
OfwZkW2X1tORmf9U9qxM8tgTHaPz/tml6O4X+S7utBNq7tOikiVbAYO2Q9XEu1phUd+2DqTxsT0L
X0jyX+qSRPk92bUilkfq6poqoKQvQN0NptLipSqqS64RhbxHT92jqrAxsApRKT5rzemKCag9j0Dj
1rdqkAeOKhy0smHitMi554ZM/u2IVCSQmKd4OqdxPXaPB1DzEUQVuR4CvJqfYz4fgbjA4sO9faaa
2AIdCmExMZtFoFkXnJypPkpzKvRtGbcVUkrycwqdGRl1dLbNvtXZzQcRVXsCUYu1lV/cj9d+132U
8JwCwD8IPQAu60bQNd5Ovr0yUy4jmfDEOQnFn7ePuPmIgsydWGTDAYaNLTX9C7gApcSUKUOrhhGS
nXbErLvdKArgEprcETX5EURcMA3mPQ3fzalPhVrUN9OfyPoBRHX0iv15D4XPFksygxo0fHPrOhvT
Ifr67uvX7xTrroxGoEVkrB7ry2XmqfL56RVFfpKO7kXnbFCJOdqUhe60pd1J4kGJicTmugx2JJ4Y
pLuF1J8rlYYKRUU5eon79i7vLl0npoqJVAV5/+EjGZxw8rnNWqDHDlxin6M2RwKWEdk7qEgUfQNM
tHnxGSAMz82AloFIAeAb3UlH7OxB3Vh7DweRkwHBOCUU8r2AaLT7NXPokzx78dqbISh8CP9Cddbd
SNzWnu1wU5j6GAQNwxiQjAuMaH8I/THs73PWmGUVWslmjy94cY5xKn6uU36HN8GdaR1mdwykrqtC
l+cawC/UFirtMqD+WKlCQGXi1w8YznEI4mPHpJLiyepSLzkoi7gkM9Aulzjx5sV5pVFb12s7/s5p
fQwm/TPkoE5Pt7PsLYCcP0x1d57/nPlDfdUl868ZMbZehFIcRB2z/bmlSIVa/BQyeQw1yhU/jkO1
YtH0Nxlcm8kRovB9uCuQP2J485yIsZxbTZL7OQje0PJjXzl2KSfweSs7dOMUATD2DM9KjXTFWItU
66iEdeQzC/L9hyG1YhfNtB2G4LEaWWFxd2nHGXCd7vdiGYwhLU1zigFhbRllN4QA5QuIcBj0gmzs
j/RClZZHIGlD//zAQf1+/2oVBDKK2EiPHak6LCqRGTF/S5ZPfBf2htQkEZ9wyFOptjkoN3+OT6tq
QfgnsbYl05izTNjDwVF/oC9qNxYsNOGDln5osSMg3PPz8mbFi1kYSnpo6IsoZ7fXarGVNjzguhob
Szp/u5nBjPCLeloMJnZTHRy35SmvMjq4Uyd9nV9I/d7d6wszzzvPMxXbK7qodWgGqU0b0bX9bzWW
QdSduXYavGODM7pr8VCbnsIx3wYdPRDHii2O+f1YZRh+dybs7VjJPHvCnQivWBOVXdcGAntlGhjs
QVgyMvRY8gE0dXxP/vBZcnHWZKA9B66mrKkqe7cbLSRiE8Fy/rEt0frm+2xrhxcsByEMFwLNuZe0
N0o5e8LHbWBYfwCo6zMV+ZXvWyadLOFiGkSFdBvgnrR/JR7eYjVBnzyxL2MtDUsmSNao4L/3nnSI
a7tNgj6IgqGWTIyxgNYWX8t5Hj+wvnXvx+PA3sjEKuwLOCaM3OecWSqpPN4dvJsJXbaaMOdh8tBz
75Gxc3t9fNrlHAQD1020qn8MBiisyRijRDHf7dVdd63KBr8etRlFTVcLq8aNcMBeG6Dbfxdyx9q3
28cuXu3XpJLemOMTvHid729gdYkWtxYDN6+ph3dZcntQSp3rP+Z//VfJmD1MJUFt1HjP522X+DNQ
9b6rB2+XNNLDkzMyqs8IE+GuqzZpIgc30bcUJkUSSQn5zMB++4rrCQktb48maordiT3nyHlMgjMy
v4fRYAO2EVnR0rIddtxK6w0zE82GcHcKVLGuhK52emJAwb0ZEG71iatTIvuTFyxdITwPoZBUJW/o
IJtnAfFf3GZ5FdX8jgXI6FLnn+bnDmnm9jdkVqrECobeSAftL7Q+SJZxjFP6SDKlVXb0Xwpzha17
faGPjvRdWgzYSg7x/jzWQBLCWd4lJLxEnY2/Egkf21IapxSfSOkFlHhvPz+I6OxO68MY32YOnvGc
IkpbQNDio+t7PrJA6Xnmdoznm5aVfCaDNxe2GCKD8B8ZsVJjHbtBNk6sbAqtPQF6ZjB9Lei/4Qvl
5xR4EfE4jKQyFsxlPmul9LyvGT/GsSiTx6wA997iwdhx4GtvIWL812DWGyOeqpJiC23FIwb3igl4
Xy2BgcNSe4vxGwoCBjXXv9gfCRQ9KgmAI5CAj86fA9TYS1Zc9kq4PylNMxNeKH/ezKp1OadiFQ12
fli448QI0Kpxp3C8Z/IpxdoXDw4KZ1k9KSQYk/H1MVWNwuV7nuVdd6eeEQHBaA/ZPI4VYzpkrX7H
ax9jrKRtHZUVQAxpoAfFLorcoZS6JD/ZCGhHOnO580IOcv3XlwhT87jBKUCveDpSaC3nxguaTpRL
I2z/Nn3AHFRN+7zh3vgbeP2k4SkyUa7dMJxM09caTTxZ+b/nNk7qCWbUEw67oJziuLYJjaAVlzKX
Ss6igra9B9O+05m3q3mw3HeLoh7wwIUlLrNypUY/ySdCvCxMQGtuunMB6eKNRimrKx7PDpu5wOC0
3MZOsfFtpyFYBJglHwr0l/OLDMDx+JB0GQyv/a4AP2l/Y0Ch+mc5n6g9GaOts0mjCsHmtuIiSw1i
Cj9OVnydfNrIwy2k2+sVL1V0D+R/aWpE6G1f8KqAuFaeltpMUFxKgeGa3ISZMx4qZfWam+8qHlV1
esEkOj5dbp39Ntjf08U0LWgOHADYd6d5o0aOUxVl3RhyfoaRCW9+EoIjrPYuAxZzuxghLwySrVWf
Fiv+ROa2OLZq5YcazMy8epyQXMrxjfSCPVwqpEddJyop9khO3ibpAdG83bX/YyfQgic1Tgh//zBf
ldVKNFCi07MIYeJL5ZFcmPlP1q0rtTGy84Co9TRjovqnGhdCCelKYeDGzQtQcbAix8jVkUQhTYAx
YkQF3kDbgYoXULIwBI6fvKsYHeVGKkD/ywh1FCwk4GTWZFI3p8yF9c6GJWBOBNr8ordHYvOfKFQ5
i29I4JixKGKLZcJki8I7crIRyNuSUc67A9iJIhQKNrCOij1ZDA8/PRMU29xv4O4+ZISandCT4LI1
ff962cUTk7NKyusXbxDvpxhKwIRzBwS0SS7DFy95Rv9YzE246w15hDwNJPv/Wmr4FqEFLkfofL8h
lVCEsjVKsNTLyZP+gBCdB8cdCdYlUl/i6umjT0afBEEboieTcs/sKUwVOUCNIS/6x4ru9SKvqZG7
l1eL+XGV6TqDYjE7bjsiHKDdicgcu5whbN5pk8h2rLgeeUPpnhy76QGj1njEBCMYUKDIIYkfkGG6
/IBL26KFwwXbhrwzH0XpS/XhZaec/0zt9/zvc4ZNX6vSceLGH6mmileAQpk1Y6loac7G0MOFTyPo
D+dt2nfa2RlKzPLQIdz5VWAlqSfl0yhZ9Fb5E3pwH5klaJ44WsnVwGJGz1Ut5mNULmuZEhdXqR+J
m/uMVBcn03ezP88CksG/iE0Fey9mU6nXCxfYoEsw3q/xOrRefofEFnI7ASwSMIdl4F1iHdiK/qvV
5CTdiAP3ShbsVoJMOthjILNuesZ3tbn1V2nrtL9kboHn2W1wTjzmgh90jcp4v4Jgq2g2RPYVQP1T
kcJU9irmHJoWxDxedF6RyZ8CPrKA3AAIo4AxUCE86TNWUE17ykzEz1bevn9Z2/gsu7nWFA82SgJ/
mFp0uB6BIc+DKqxZqAZw1Bio9raqwibJAktK83TgksKD7V6+V7nJ/yTnrTJ59k+v/b+rsOl8F9XT
YlSIUG/aZbJLVHnEJD1vXq1IMVYCebwSRLdqclIjWmMcdPVZYVcPn0qGSlypc9YsIFjmGjZE1oPI
Ao4ovIViAWVn2vJnwDeohuNUzWkkS7A7PdEu9nmbrXyPtGXubuL63p8WjDFacNQ2nn6aZUJCq775
Y3Jy5rg/FWtrma2ALeLGJl9z0FuXA5wyNsuPgUEYK/grTdtbnYwktg92isDfabaXdOOV3L6qoLCL
LMEdk+vE6MODbMBPg3DnhpdnzrF5Vxe3V8JoNr6LQ0a563ltI+ZaeL57q7TrY3MF0ReKokpTkXGX
Yo4JhydF/x/zHvZTERDC716mm9oZmZjgIyXDPsXB0tz9FvhJIMSICUlTpYt3RQklFCPsnbXkgwuz
ytwqFGv6FGcOT9V9KiANjiwNBD5UObuLm3AeDyhfItUqAcr/5fTsWYqQXUuw7urWX7+Z7cJqv3VY
DdXTXIDamE7/R3JQF/1TEtNEv7mRv4BbBIuH4bdeRoUmJq+vj391zAI9GGHJmL+aJVlbefGcvCC7
22DjIxkevtqiU27EhqDdgYn1SGJpl11gUXXKWBjrwNArwvBUEoJ56bOD2Mx+I2RgovFYAhTdlnzU
KkNp7PkDvtMHVSGCV0td2xJQxuIMLgLN1BnC4HctfuE+is3xm3HgkkfhZVIOkGqDAz84EQ02mUl0
UNThQS3ax3VlJnrRddcVUe/+rqSoQ9o29JoxtF6BS8DCSDi9FFBifadWNngog0gQmjB22fNigqih
qLU5yl6xmPYvnxx/L6BVXph0kgQsmyI3PplI12YQm0s1gND+UgPxWIcnOAxGS17UM4psAg0GFPax
bQdaBGNu20qJToWY20ezCcQxoATuw/2SVU97Dj7SOjlWuaHX6vy5Io9VFWdblj7j3G3WFVqhgM/l
iOOz4W1ucCgf3S38dUsx7fgMtsqVFCLtAQSpZPDwnQHwEQab3qwgWM6Nahe8pCXp22yMCdjT+oK9
cYj2btv+fAWLgIu9xmpJjPiFrRYueGq368i/ExT+XMF7290ljssfg+or6rqZDYKVRZNp7PWC2Mfr
NOJM4XpktS6I44dmy0Ll8an++Hi2f7t8eJTiduQ8BzgqOVlZWW504u5RB+W3pE2azj/tdDtWHJKa
+yj5npX4VtWlQU0cZ/cra+52+FChDr4OhEaYoDOxo9Y5FBkP1f+4RiB0409RLJrlLwgXJVKMaW2Q
WN/ejiBPL6A/j+ESUwEG1/ieeU+kGbsnMTSleKaL0DglTTzDlp062OLCxWRXJTs01wd1nOi/ZZ4W
502jXthP1oGh7TZhHd8b5b/46K0GttzdI2F54HU8vav8eg2392Ek+bJt+icCCAn5bTD4Wk8C+Fnt
qiECr/tNJEuYJmy5FL+J3MeTIIgV2QY9cAfJ5nqFV8yFeKGm2rch4CnNtis4z9ze2CKVMeH3V8JS
A6716vEHvuQeHXfrv74AuFhkIyYTxYFCBei262rE3nVGtGPl4jo4VtBv/l2B09OD+DgvCoQ6WRxP
F4p/I4bj9YsXcl88ZgEGXxSFaMwhuCBwaTdMUVfZdc9Ia9k+O5tOBE7mu9xGMc1S3CVZzp8uh44S
1MrJgYZrl0iFjU3quFsm5c/0z2hDeg7lNQm8HrCPcgFi5YaaXEPdRcgHBqViL8RpeaWZrZ4Xj+lp
eFJ39M72yZrDkvFaoSnHYPvrrMX1wQFHLgDg0sa0xOoHBJiPQWxYgTv3p3WbzcIjX5bXrS9hjLQT
a3Oa/qA19QMZcixhyG9t9Zhep72U9cUhmb6wzM5H5YI2T87ymZL1UkxTN6LEHK74dOre/aCoGW5U
oNRGbAKH4/boECGI1HuRGruOhGdRHOMQXK55laNe+gQBvmoyYrypKk9yuSpwJNPYYWc69EAk1rPf
pytYI+0b5xIAoi+IMujWZAI0udm+DwcBU7LAlxRXpLkBc1ZAKvLCfaHx1xqkMRBXrwbNOfhNa5F0
qq7mcjc5tQbCEya0G9x3fq9ujh+5ZMN50l3JgDcFE5AXUQnL9+FrnqlTrqIlLkIFwuWx90ZoYemp
65IB5DsFcaII/xR9xJKJrecX7m73ZMpJRGwj6A5Wex058lqYHm2YJ8WcLQZgawqOh7Qhs+nrIvaz
XzEgL2yxzp8z6DIDVa+Qq+YXK2lLDB6kQm8VECzv9GgkmHU/CxMWUTJHgmnC/cKGZLiQepK68V9v
g4jUDbg3RgHPiy4ahIFWcDGJNsq2/bdwSouuYHO9P5BqGVAWarjivjj3gHsIWc9Pu0zkFNGIA8na
fDC1NvP4jpqPfrVCDpvQbILdTco8XIvgBRJ/QRwcBMJB9VJDOIcPEtLdxT632dBJrTOYNvdahIDh
z8r60y7H7EvvhrECsUyZPsLCE3exDn6OWIQLS8Yzf1ytROEs5vEl8KbI/+4rOdlS9z/m6B+1LVam
tAmyLJy5Zn5UsZ6FeY2Ssge/+Ea9xWs/8kHjNm8QKtSeq/idDTqgQY9aYq0m2V5ih1NssYaaq2Jv
JdvAnJTTYtfW54TsSC008Njv8+R1w6lxwtvzsPtHsAKqmpepwbkN1GLE+e4uHrsTOkqYLLVemyM3
k3aVfsF5u8fEFjH40P5Wn3ZRHf8ELkvaFvytd9wIyujlnMoyxo5IM/Sve3lMvkgyVZRi5QxitSUc
HUxbTKCSVvDWhlKyEApR8mDvkqjfzQ3U5G5R5iknQ87jzeZ8nl1y/mhMPg1xAlmVTjJnPTiVHTbP
YJvXfNYAGjHZCGtKXIO8YcJZhwkrYHrRdBRsoI1bpK/FESMjaMOKtS4kJ0ff7rpQUXawIk0ceiHI
kfnrftwfx7+jWVe4vzeZtyNgOBkztUokxMO1/OVWzT5UlfU2mLZaeY/KpPTUXN71yf1zTeSAPJua
0AjOIycg7+j9uZuXdG24gDIClu16HXIexujFIRPOfwd969y5qUVSrXyY0zAf3jqbB6r3h0VU5whZ
dnXxECplSQs39VSD9CGN0X2B9fvTggQw4kFhrUzuW02CTtLZBajUjDF4DO6ftJTthsHEqaSBy77z
1NSxzGqwY9I5VI+jKSIK/tqCMI1oKBNgx+rOGBXoy0pEQhhy8c4TiEBN3MnSCb+Qr2k8pTGDC7Ts
bgn+7yQVhJa1aLNbFafxTb+Ye5YWreeC/ZONz+x/TrM3dVlr667FXB1e2fwlOpQ1KXmLQBgp/APP
b9c6rP95GtUDYOKreqjc4v16KaD9yBuKIwUmu8l5V1lhlev/XJk+yMBZVyVw9oKlRa20waN/LbET
oLt0fz1PsqXm+ATZyUd74cVYBmiL64oJImkh83mv8KkGSESb35NPtePDfyq40fEIwKyCcUESSaxF
Q9HO4dj2ME3jiG3jAetkvfBlFhOiv55xf6/7/+wlmD2sXQu9AVhXQltHAqiQCP2oTo87qd9VwIAj
eSJkRZZi5JHuNuAI7r12Jf8prGoDvwhptEyPBht9BuiPLyugm3aLsH0qdaaibbn/Lstklu6m8xl7
694O0/N4zwvvYpn5RMux6T9axE0VhqBz+zIuBRuumXenQpBRLaoFhIMwLZSlEtjrAPQ+KOt12u0q
c++B5ojo81rrf0Ez8y2hLU3xNpuZfEXy9S2TLprc0bd2jkRWkvnKBhjzcYXYPNL2jX6IsNG4trW7
l9AIXCie4gDY4EOO6eHKt/USqGKvdbM8p0TvXiqFxvsXZYUXgl3ebzoqVTj+ulk7MtEIUU9IvNGU
0gQzJdaKcYWPcSv5Enu897lOl9ulGrLhdrsMkOqlb9YoHcslpYLInHfkcatXwY0xPYjEb2MjIL8C
gXSZ8dLV6jKNh0eEboIkH1pKACUlBq+BwBtr746uc6FgVFZpJJiDnZpq5HUsMdFrHxgI2+ZTuBK1
uw9QsK/mguHTE5sDwUQDMJdinG3ln8uISkKwCS2N5QHhKWlhylj7wwHnsGoJ2DUqh0JZt4THOBN3
rPmSK63H/a8eld9czogo6EAszRN4AUQMAsz8Wl4vWR8E2zmWdjNtYwCa0BOMp/U9LgK9iOIA2+Ll
U6k6M5HAAuhCIOXmUyT6ErVR1Q6ANwl2G+85bDQm8EtCjPV6RL4iQa/oZ+OPlSKT5nh/y3uaRArL
fjkzhwikXNtYhVq8SN3DsBaRplAHL16fYdr1fs6xLP3hahffO7ek0QWnc/vv9xTy9NTv7LXkzlCb
+ZKxm+L0tPVbfsO2fcfNgBG3reQBHmiccYPUMk80n63PGnzmWe1qjzRM/Mowk2fzgc8QJOsabHHS
kuI7e7GBz4tEh7Nk3o3qOea9SZHGAtb+wTRM13SvkA6vGxM/7VIXKsVbjrPxaknkdvlu7woD26ec
HXXZp9KaYILXDHCUZV9jaYY/2Ycl8OAR5Ondkn8jpnpOr/D8lLFPIpnkbOaWm/7xqu67+A3tlJuf
aDKC8Xdd+UiCzzCvXpcg8vyoNf2qvF1O37e9cvC0pLWH2ajWXBeep0csO/i8ZCG+KbkhRXP0phPO
mD9Yx8hLtlQllSB5RKU5v4AnOiedTLx3wFtgube+JCzq4mwbgLHpVFhqX+WxZCazUNy64OCr9NoK
WMvbNEBq0oIk4E+Sv6X4B0sXNEhkm7A6lmq2LKcUqp+MjGdTEM9IbkZD+XCMkLPQ4c3q11nge1f1
gjui+3gbHs/tzQmlrt9BMxQujRY/3x/JMfJoH5r2YJ/yDyY5r+8f53ygKbKwYbumNeBUNiWAaAwT
WwC18/D+VCXH3XkXk6V9rd9h3/Uskaklhmj8nBJAehzWwRSnGdQskN2b7wZq/+Oml7XQoqvpeagT
nPLuNdmsr0d33d860EhuY1OEiRemaxKsewbwSeRD1Pf1FYGYX7VsjkdK0QSbYtUbujh4/jefb6P1
XWEPcZzYmKWMQESrPVc9ugchdV3vk342yxNbd4yd7w/MDkNwzgDeJoOytmCoXHYjySJop3bBTwgj
89jHysM0Kt14qu4TlkabgIII/tUi12o9LZGM9ceDK5ubRXLPH3neM8ixO64YWopOca6FGjPNR80R
sv8Xepgpa9wQGT7itNy4UPqs6SPJDscCy289DI1iAuPVYzFmV0NgIP0CkJbr86yocdwnb29ZLNk+
pdgt53s5jT2CIeZg70EGf/crQ1m7w2RFtSB2YDp67BGiwsk0Y2SukoOeOf0hH+w129sB4FoN8Ep1
ws/wYoR16xGSisj78auBlqXI6ZIUGfWcRoYKL/O4BHXWzRnTSNH20ymF0NBLQQoJkzNAJeKeOrr5
DoALVJfXUMU+flg0+6C1FzqUdEVcq9+asZlLHwMV0XYhWaIpCYMu3qF8bXID+HYo1OwmlEZEcNYU
6xasDe8Qh/MX9YEh7GNlOZDq3KGPOE5fEqoQp7f1/BA90guKyUF749PgBXOxEqmqitN0L9sazz8J
M+Oqj7qbv+K5NS3Q99rkZg/U8eT4hb/X83I2QmzCeQvwlCiy8H0GBSW7sI7RFbsGFXtadGTbrMyU
nXnYMBWz+hDY/DQemxji9LNWkpeEwSFQBqaL354M+DTc9/aKaN6uXCwQVfLzZeQCWdGOZZ8ogtFw
R+WxLPK7I3dEvM3jCxiS4v5r8aMWqQhCBEEMmHNa40BNe+w1Fw5bOg+6EYvZ8rdaBv/3vBDPXlNB
cx6FjS/1sfI/loYESEvRY2jIpHGht236p3ku1FQOxhgobLqUNvsgmFTsRanJUV5NfrVN21b2sMpu
EE6J9ak6JxhxWDh/rDfegUBZNJRNwbSJWoHUVlUy6H1IcXLmu4VWpjVo1WjVQWFBfR49vqGXkFQU
j+aoQzmXrdv4GRTO7EZauDTYC+Wk088+4+6e9Lfl4WIqMbusG+QGWYHIAZTMATxbW3jNtyAKHgLL
vR14p8wX2SlDQPlbBZFv46t36vcBwSATXNqGLzhHiF6JFyU7NURTy1/JgBRIwCBMe+hw/9mUSlrh
awNZLK8YnfvtVNfYoXBZMRRINMBPBH3wTskj5uyrnRpwdt7N3o+In5SW1Y7o+KQrd5rbrgKutiTD
5ItRE+6QNZifqrhnJisKFG+SO/d8eDrWZ3mJgcXSUjZ3HKs1senyxHYkAgOH5uDdnUgQs3bK7zlk
So8Pw8g2/+j01jslaboOW5+0eBF/CcRn8DY4HP1ST2TE3okiZQv1uoMymYFlrdh3/DIEFzHQV6Nd
7T22puUW9K+tImQbN/vGSMNZmYHJWSgyByXbY0ZMvA6Tt+vA1CkeXxSUk/toWb79srgVSmFoII3J
xwGkz0qLE0mEs2TlGjSN7UIuFjBagswfigfrM65UjqOylmnsx3hRaduZkEbOqPAU5yp2WMF4A7NR
8T5t7r2uUGbvd/gg7Y8yt+ulB2lKq/v3U7Q6G+BxouX/IR4z3atKoDiJmmfn9cs0iYyMu2faqdHN
KVCPJ5diPH+bRAkNyDA09o2SfZ/DiemMOfVPoSDxmEjTOSQPzfMwZnoph3bj4/R3GeRg2N22zWQX
2lzbvYvYNzD6tfuWXQ+IVc+rXbRMZbeGMXO+j3EMb3/3hrLnDZQnL+/0wYv/BDVu9V1yYFHWTVEs
RmRcvuxcOsyX/m/DN7qcE2WjvmeJDdcTLJUZle9ssIgCOiQbOCe8e0avGFJHZD9rlepjzx5xy7xc
gbZBIaHTzRYZSdYYDNmdEBJY3tJCIQ7W0rdTKrkbTPbyqmoSJTzMvkE4oXox3b38J2NSVAMyZIFT
VQ5jcb3Y+FRGDPW/kQE4ndtgF6tJ/oCSQ+I5ciIfITLHY/PQ/0D5nfTyZqBo4ooD06f4gkcobk4k
KbxJ8LAb7B3QSicoXH9IbXUG6gxTofJXS6jsuG2UdR0/yxLUtbF7C21UH66SLxdIu3rMMlLfbASw
3am7HN1a4xV3Is81KkL1Rrh+IyCnn2ClMI9Cf4AKRkhnVHRLBQ5uSdZyVGOjfXJnl5ovSLciS4Mr
70GGuVBggkK7u0R+JRrEmed60xUmAUYxmhQ6MWnr9oiOYWW4tR96u4ZLIGbRdTMSbZ/KBlwigGcz
FoQk7Ou4Ccm3dJ3rAvgBJyoZ9NX7llJcsTWjuezc+djKevmk+fWhoTTyx1xT9fsERr+y7ptb+F2c
bJfD1j47ii3jpZciIrK/YvvTSbXvmmfh77dzw9glDW0PQWKhlMD/IHVzjr7MnGywq6Tp61gSkr3B
auh+GASvjfqSCKSEBRkgQbmZjKNEY+KdDwZbDxRl6lv141VH43j1SfPDhdFwMtkPoPauVCU2b8t8
s9/+SCciDo+jS1Zd/D0YMbZe4pPUvA5d4fzJMbsno2fe6V5CPTUHdNGrerTdARwzEbqJOY/rq7yV
NL5hgoCrMX9eQPt9Gy3XgcyvJp+TFcUPR9aIVHCjzdIttbxU2zMujac/MsDR4PKHHTpM6OysxjRI
P3Dp2bvdJtQ7W4MQkkVVvJyjdd72ceVDg0l8J2POoUgw9FxuG2jffgUcdVOHxwoZaD/g7o0lBnjh
k/EaZb3zPKW+kyd6SvtO+c+CoHAO6LHLKtLd538U1YgAvPYfdEG11uolWsDVX+z8tPbsjCIhTFdy
99QO8RGYvSo90mQWEZGSP+1D+UYHq2oj0fQYnu4XVO6ZWcWkCiQ1fTaP6fatGzvOqkM/SuII60YN
vVDy0N/7727TAO8mBLu6Yb/nW58P7DTo38kn+2XKBuochPc0OKxri8As0Sq6SHpVr+pFYHuR6VfP
4ht/i+4MoEBtieBhFRy/636igxaqoEpSP3LD32Bzu9BujthY52leh5Eq43s31uFjLa2Iol8ic03u
HyaTKDHSIlcXRQ4dYLEFs/bFSQC9r++vipULXYGej/LjR3HaeoWn0rxFNbZZF1P6RErsbVO4gFos
0PLgs+XTKT3Y97VAsTkJcOdBsjPODXEihCPQRbrzctdHtSiyrvI4T65hEg7Qmm0W1Y3cPl+1msPh
Hzd+YZBa57X/XD8n/Fr3HoAlhP7A/kUyRVqYKegQwiUhzTYUwkVKkJ7OU4eAHMPC8qJNQpFBNGtu
Ow0p4kSrQPTMtrzyv5qRAgBG2NNlhTjUbjwvFG0Lcbqev1xGJIg4YzheZrzq9NDhvA9kGkbW8BDb
nDyjDxHDDo5KI4TitFVgDsGs73IHpe1iZHVDpYJ5hK3maGaLC/M80rzQgo2eO850c8n1zQ+S6aD0
esFcY+lXIdN+r3iM82VMUj8A3lw/FODoi7SFv4+giafufZndcsqCPdi1RsToON0aPCiOygCRagKe
ULv8D2fXNRCGaf+wZK41yUzExmhYAUiM5h57CbW7kdpRhtCZMtdl+BQxSQKhP47ikJDoS8oBmFHc
PGajrp/bNKMKxY9NKzfZfytr1B0pkIEKvfDd3hQBkC1x65kOYG+j8m8elcGuoPEp3z49o0ZS6KpN
s9o5C56VHVhnk8nSRY/mUAFOlQCItAqvMW5bLaFm7DThj2yhYIC8NaFd2wu+9lo5XUyPcxiifcw3
6UmVQpCrYEm+6Vg+n/hkpWte9HzeneWIfHleF51Tcz7bx2CJERw9ofskAuounvzsWy3lcH2VyxSN
edn51X88L93vDhawzDTw8zJV3I5AdYjWzfYPrO6BmTTpd8OMAH/wNMg0Ldi25MCyIQzw0VhrtpaT
/Djygiy3I6wYY+SQOZ2Q5IrySgGZkT95Oect9GMRdSeDup5/7Lbp8JzChsGcYbo4cSSPDZ7JHvN9
MiPjD3GL9toqVgdChATHM3L7y5aBMNAs5FHUrKMV9oaGwbv+R2JFKkQT71415YFxybamoReryeFy
vK8mEw3+yvbRGlXixTrAszYHDEFzvdBSzilRhHUsXRTQU1kq8hThzM0Br4sHoEcWrNl6vOgt1Y/X
pjmR7h94d8a7EN074/zah7DQ8et+khJi1vJHCsy1ywwuj3dy7pDxP10s4Tuco1pF2w9pU3ahuTEp
OS9iFjPYg4Xace/v990dndBFrXB6STSwZAsZIKf9h+zAHeHRvtnpcOp723gMxRFvcvJhFeYHn8OE
1/KsJjJjEa4dhpGYhvClV9Xen0iAHQ7ltZnFvI0KegJ6FdhP3hl8Pdnj0RKp83/4dAUBkLRjICec
3K+yXjabMDFj1jhfs++4PnNmVDo3yeLV2SzClGpwiTp25SSAKsxo6WGtU2YW7dg2FmNXIyG21rSf
uEO3i8P0CHdfGxC6F7Pn0+qKgmE8vEPCvdQTJnWSRvtVehK5Xu3SZfYcPROxdhaEIjeOrfQI2WkT
WGEJVG3PUHoehdEQF6eNvpEBJzK5zqmkoQU8VgJSGappXiHmH4IX01g+wxy4+PRb1fhMqcvlCcVv
8CctFb5Aj6g+eVgBcey6h4JP/xpF7aRma2w2fKtq+15BpGFqyWnlXsvSEO4ekh8QJOWjLPdl3ZQM
4RhiSzJSOJfLUwgf/mgDUcSH/+LITTtd77vRkGBxh0ljlz95V2yZFNDt+6ToTNrkU4jaohCbxF5J
vjwa7PRt4VuweeMw9bP3h9R8bad1fG9ab+Hh0+2K1YQTsPDInsJqsNLN5IDE9Eyp/AqRj10ytO8Y
fyxpheoRGPIohETGFfWcTv4GGt9Tfy1e+IJ46xOr7kTc8Jt00y+9gjk66ZyxfecNMrdw8p0ZbNu0
+vNCHuVauy0MhO7vS1GRMYFdVB9IXbexK93+lCNBQQqvqv42JnWueqiI8EnnxHTp2HGLNdZDCOPy
jmYichN46vw1blK0pDe15sSkqOjn47stksuVnikrD1Vu6sw5JUEywM9j68+bMc8c4TxZHai28BAx
ka+qflaSpOFXW7A8LoCFJJcxn6YoO+6euWz13+21Op8LZSp8dL6vnepD48iPDc5SfaZ1cF+pyazC
N/uYcOpGtJLzPPDFLMkoM3yd0I6DJE+6wBiPKflPIpwbxqw+HmR+kBxxYPkqluYh1ANnAVNnfb85
IZV04xcrd/AlGMR0GCzBdDeWoyYnZ7OzFGXGxcGn88beXWBwrkfbnzlGNUe+LftD560BGbiKekY1
VwZRFiWXHrF4onuv11ywXM0cH65QKEqks+X494pPfUUiVzUTIIbdbL1+cHHQzoUnXWALuo1BVQW6
rDFER3kqKEc8/8eZAJhrbsR46Ng9fYqvmx/QrUWZNENcaUKwz/KglovjuuuRC3fSzGK5T1WEMWoj
MIf3u2I4lPG28NrCTGnVcsus/nfJQKFo8qNgivzwnh9okv9Ll4vhNFencajet5Pcs5ivZgzd9N3B
4uDB9DnDySeosoS0QebBd8oshtWcFQMIFjZEdATJisES9Cseas8YDUe4bGQdGduU3pv6Jcm5ZTmp
aNV6p0YRvUBfsFIPw0Lf3r3z8Th+sZucuokrtK1jHaknwpnKnilm4nnu5PzECt3rAR2fsXHUnLck
aRoAMvB4Bicomjk8jMh/tTlFLSiyMXzrcmjkh8PT2LnE2c79kx4QMBLOVxbD4hWoF1L70jRLlsbN
nw+vFrjHUFL6kLfKcc7m2UmA26yLuNopxRWwhxFk/gtPX9SiZmlqhfwrrmUbBGG6x7Q/pnkemAxR
Rg7IHzRZ1CfhRhKuMng5OCQD/V8xcdIDZ9cOWKJM3zkWK+0s6feys6ReEObCH0oNcuv+1q5yk0U5
7Q3Xj3pTkEwJvn1TvDWmb/VuvUtFQiHxoE1xnJnXt6Xqjwkefgzv1W/8ZuddVoZoVvraZRrePOfU
8EDDWV7LFvHnVVgUyBP4ThGsTFSk5Si29bbhrvp3kCtjc8f7hMHPZXDtWEp6OasbPCB1mDNjzcQH
kX3YUx7HhSYswa5a/vSgl6Koo1b5DFAZRETZAb1BTyluPdB6JYU4oETD+/UoiDHaJg6GX1Un+j+f
u7AVt9Ib0zf1wvV9cQ+qFdCC68hPv7h94vv2gJxqCcncmdSs7vqaWZDHUvU159Q2XevDq/l50irD
ENF/Zc1vUMAkUidal/ILQKs5TH6ftZq8GAtApj7BUmyJEWb5DchBNfsNqE5RqHPKp07BWxC6Z4Jh
BTs25jhiBl2UGh2YpHqGMGuGo9FeqUQB9mBruiGoxueIfGBAk2VNNWcC5VDjx/NRk7GE/JYl669I
dNymJfHunfoKJeAlW0dDeODOJ+uFU3Ee6/MufKYEwHdz6qcPyNmkyByk9h+rqavPm+C0V6w+cQ6f
Lo2kRRrhOD+hwBLZxDoRbhW55UOXoowEcM9q7t5CKotWE4aIAsbI718qYnO5IbsW4j1ECKqk2BvD
E7FfNTLMBcmcx73mY1EUOqUZD3ZBduztYLmHtVudJhik0aozM/95I2WuauH6aTrchsXmIMSTE9kK
56vglXgRYMh3Aw2yHdkJUzGlS37STjK6AFSnlxCzzWT/cT4gQwA5ytyTm1Zji5yI8FMT+ThtzYzJ
+ecSU71iK2VO/j7HKeUzBMfaevK1spJg5oGwiM+7E3aErlbzDq4wX5Pcbf3SJugTsFGj+xTk/ohH
PTqeAuuczkJ+Aznb/fN/4mlb7DSFBamA/4hrB1qqh9vFvIxVSaY0FLnHWxgSg7uMf42gNeag47IV
+Gm2+FarcfTYbtrJr7dhC+sMg9Fr7LDIBFGL9szrkx5UKpw3uVAR5YFUSz89dI32Zut3UXbFyiTb
5oApxRP01UccpNpiiKVSFpXdsaoaP1hb8ycgbNFOjm8oIqcb19yvBl1+yjJsFzSFUL5NHfdcbASB
QD3mPWC+xA0Yd97xB4HhtrbnaU4lHCPSn9rYKrNcjcTmLK8Etj0rQzeYoyH7aFSM+Azu2v+7q5nJ
WRISqYG9rvebIJRGwBwShEUVdjuzOnIeKXd6Z8MPr1lnGSL/gZg2V7Rbw1prBhTfsOzOKjLJTkBX
VGpnOIAzWu8mr6K4m993Hyt3lzh17KctXEv3nVcpBkk0b8UPMUprC3dILYnYplTWXke88t+kIZ0O
RTEOxTO2KJ9DkmNKGHB6HD30iSE+AiqFACKS2p8/RThybwv5iE1SJgGQnUn4jeSKOh1RKpshZgyT
JDSBvzNQWxBHa9BRqd4/EDQSwlEboXS0P6UtqKvzqaeCm/xjUnd6QZJl/01vLY8uKe8ZoH2XZ/VF
OJxILO0A+4xaQ84YgSxt/B4gt/GTiAXO/jmS1uE46Feem4VvqY/XFtP0mPjDnujgaNxDf+QKl70u
SnY7lbi78Hw4H9TQoZjVwVW5FkpF0vLPGwZnUwc/Qcisz+BYc/PxTRpMgkntPIXKhelkGEMKWoEt
xUiaUWf1AHxslQ8HbLrNY+qSeC9gheLIN8fKs3XreKkOxYMV8GYvnykVdSJzWmRVqVYZYlF5eefI
TNbIzxxTrVRfxvn1z9X/Pa1vS9yO1qwCuVOfId1BqmSXlS6i9cuG02Tbc2Q31r63NzKIuqzLC2WW
946rpuzbH4MFuZbXvA2NMoEP354Q6OhU4UdD2008CBy+01vVQ9AAPMRWjU467dR09Nfkx+5gdcHr
GBV9CRu8+f8UiA5DyG8Oqhk4iNkk8x/6lfPF0yKHTmALnUf5g6H8cg7hHPA4rizBWn5eRGj1L2jw
jWfa6j7fd83np6c+QIQAfNS8vQ2IEp5qWWk//fFk9S207w5gBvZMCGvLHsfOWkgenReAHfD08Ptc
hjCjlmCfG0ORxMFybOAakxVand6hTWhtmZuikE5x5Kkf0yueyK6voK+IfaoKf7OALKFCzzjAN+9K
41MVwEVkF3QnCLNtIyXds5ysPnrTgupCgFfPZlj4GFjJB94LdT4vZ2LOq1b/BDQrgO56I4fKLM7K
RtWnm8wvaEY5HRjbf4APHpcm6wjQsIbspC/t68aLGd3Nv0s+rVhfMb6C+7cx7AN0HeWC97453f57
2BUDN2tWbkrhe8UCzFG2TcQMhDxV/v0FwsYFg600+8P3FleHueujx1jaXE3NX5cdsDRislF6t7TE
pZ6S4TF9TEb9R+uUonzCRgwhQgCbLFbqC+r+Id3heQ5SJ2PdEci8waIgjpZdOaWfy1L8X6a8RRuq
2p/ey+45Gwg8GjZRBzZzU35M9HoxBbIjnc4HeiiYSASFDJfmmmGjpmLvOJnNnrur7yyLViDhMgtO
sakBnLmMTtQFSsvMhyjJxktnTQJal4WZT5DKNLz29BxyvIHDJKjOTmjsKtVF2fckEcES1wfqw4Tr
yAv28Jv7oaOA308ptHzryfGjZnp4XttY6mVsYrWNJCJOjbYL3fQ1TK/1bbfoKA/zCtZScWRF2USH
h4d74m4v+oUdvm2EuVxC5gYtsMOUQEtLxe11iI35p+YpCfHvK+NCK7RVTohGpyvUMT/1/mMiiAAl
QeFjCGWazUFxTm48QekmD8f3puit1nxPd8njbqBbT6Oo+o5IAVFWw3UxagEUH/UCwQR94qi1yPkI
eWFKB8ks6/WqX0uXSV6iC4QVrbJ2lPpfWCv2khHpoKsPACnpclGDIEwO7vuF/ghK7ncNozz7I41m
8OSB9pRXQswaPfP0d0B97mlcpe0cJGd2PMJIfA5bm/i/6Tre5O4/GM4ZKCkh05oSkbUDJI7aECn5
LUMPViTf1ONQU6q8hbKQAN90ZZfyAoMHdFkslPnTiXYA90S+bP2TVQtLItfOkA1PHnnBx5VbKmnp
0Uppxi22BGxi+ntLLAgUrEMw0pwpfzIOzQcCZ43XBEA3URlOwiOdvPXAua+YlZUTXRU68TNveseu
4lO6tdsM4PCVR6Q4nFSoA08Kc5FGsyqWlN8R0FjyVqvZu9dwfOBgf6DnFnDLFmB1oV2Ed9FkKGEe
a2Y1qV2SrrY6PAoVYEHY6HCWP7G7cx7cX/flOg2TI2ALvbUtlwfk6jQLIDtwh5S/rH5vz/PyshHE
ApTsn+3XcPZDXIun06MdasBBYcOgy32RwpQkz8tHDeI/5Mt/eaKRSZfpDehQN/g8aY9BDDJEcfoz
3CyLypnniu/yhY5yA6hzyojC5UOIewnM4z0MWZ7ymvFG41KEIHlPF533qVNwFmv/CV8smvjcSgHA
/Jh18r9N34g2Alha0ptpw/hivyMloikHJ5eo3goZqrkHHV5S0dNkz0w8IPn93iacNgA9EU9/Uj8y
HDVAsM1py3k2IRIRx8CEmr1QLuDRKfyZ2+EH654mKAizX3nkV8xJNjTwDVDXNkD19xZn98cpAwWt
msEPFezysHVrGXH5j5Kl60//Ve5bpYOrg97BHamhTzGjelfNK4HkKKSzdr/PgjG22MklUzKzcjcs
9HSH8RkdqKSG2CL646+GshYYYZDOfN+t6chFth16fP4ks9SqJkZSXJOXmIsagq8ehnsuJHdmDb11
+XAVK8YCVT1CsSBNVSuSFvMF8qWEilQMHF6Xf6dh5ZN3zgbL7QDAyjH18IRPfisa5TN17UB0NuIU
OYs16gUCnz8sYkAjl2UxtRKgpBsYKy7hUapUOEsJZm+AEZOCIGaHgc9WJXlISesBMutK2hjDyMhI
hjOcd94jBdsVboJ58yHvNzSNFl7WRZCqfvlmKIYI31dbekpy+fTqpdVzsC9t+q2jmA0cbrlSyixf
flhHbxrwTgc0BNNRZ+MZB1JFNuC3TcHxG7J+8mpqXiH04L3UyGLHuSXSae97UtaeKsRD96tVap6V
ipPqj7sQq/aOSlTCpYPmdjoYF+RfxlmV/8X3+jL1J2uHiAUKRu5APVaegLyPkA6A8UnVl4UMKMvi
VUZHliehsiAjGln0dMheHkgPZOpd1+uWmZxHJ+sLa5dXiiVFKPlxpfUKIpGuxpPbcu7bOBgqfcGl
F46eun/yEkc4wLZLCXfZz0Bz6cKJVYuwwNGTTu7C5fkDmm0KDud88RZjeY7AW0AUvklVGfce9rXX
WkWPYlU6u4M/QJYGBI//5E539tdgG5VaFI0mxKqNEXDjZWEyJDJxvSs/gn1D8cCvev/giiT+wh01
mGSwC/QjwM9sXzNDpVCnmhnqMZLc4WAtUFLjF5HPvoy+Xg3rOwMD+8k6OdTIsA2qjJu1op+O4P6+
8G4+extBqKNdwaULvsQcToVr5wX1klZTzHNbA7kwOGSlHuHvLk26Irjx/YR+G9JYx2bE0ljf4kVg
F1f77z2yt1zFxCqWIcBjwGIsFVabrVLwCBKSDj8+24iN6GZ8GfSp2F7AlUBqrnvf5QE5gs3P21On
+C4xCAcGbh3Wb6UiecjnJ5LbfRRrkixA/z3+aAZcDXKBS6uunVkISfc+1NQ/HtOwd9fXs/+mYhFj
NXlAlH0uX5vnr2zSRo5h9NHEFHXwF2h+velx8po/ksDdyjJoFpVU1n0oVhQvdXr+ENc4iYj+wzld
5ICfi5sa8UKK6pqZ2GhMRPwMCjYcyJvsHFV/VdUvh9/ZvgZIZnSZkvtMcNTIICn3oY56oy52eld3
ROwrGvbqRtidaOoZs/3u1TVAr+4rlK8krfGD0t8/fVSYkGHj4QElS5oMJU2Z9gGbXyuTXZ7+R1+j
jwRTb/3BuKBTZG0VtX/caOXIFEl1b45SqQ+ROPVoIq+uZe9C7Y7svx8ZYYVhTMbnaA50Pa0Pdroh
sb0GtPSJZSYzZbfMOZZGj+Qb0uKdbGHEWcUNaM284d9wF4MeX8JuwTVPX+wivjXpuN1LRZlljYXp
hzjm3QrYGxaprppE95gGpaHfVC63WnqXz4MfS1HLX14+G9UAM6cZExhu96Ly3NpeWBKUY/TnZRJV
UO86yckC6gx9hzxkTvDiFLea4e6MKNC0PlKdmkhJiy4hvUX1S7JV0/BoHj/mPuy0kf/Yo+SfWrgw
/AwJtP6BOPSMcCWyiOmPnODuQivxBKhJRbmocoa1K+XnrgfiTWC3yfC51VCnKvGp0e4yt3dbaRsj
y0zJBrhIuFwl4EeHigRtZNLj2ue05Zqaqd09FHmwoGZxS95ASn3QmFW87MjoCiTI6p27jwT470x8
yLQ0oQLIO+J3/nkMOXLR6N8G9N6jJR1z5azzb207YTLxs5mBEBmfyv97t9wbmC/uBFKYkHs/ukXX
2xyahZ8h7Bd7JR5FAfhh6GSnts8CgzZcyIaZz0Q5Nis8o5FZgTLKTduWMkOEBqPj6NX+ZN+4TVNt
Jd/tpORuAw7bydC5o8/6fJULydZRpg5Lq1C+LlSHaBEbgUHYrJc48+nWo/zuHGvGpAspCPTo1MnA
fVICVd9rs0uZorcFH3Fk5ARKyvJiV1WbLZurwzhEHYlHLXvqcqOD0b71LfjUGFlmKlc9Nh43NzdO
gmC4g+Pv72LV0RHqBhWuc2NC1izaH0tnP5VOTpe9XB5OiTiPOY/JKwxZJp2bPirW1b47kVQVJA6n
45nQGCu0PVtHQj3qimQHCzBJ6WLyGBVKZmdoKx2NjgC7gs1dUoy8bKf/UkcvUVWs705dCq5lFxKu
6TsTHp3IM+onGpduWtOtI9Lnjwf3+1w/QHv/qB8UUv7UX0/lTlMGMW7FfFOwOBkwk7qTpliTvse5
rR2M3kpm+aX2BMIAafo2EWd0m4JruvQqa61MMwdhyRKTeSGjZNjFRW8VnIMaOxqECEL3JW+mD8pA
mjl1hzDuMSCV7PBZvEGKrWEK9G8Rp8MrssvBD04gJqMeWbQ8F7BpbaSVDVvvcxjcKj3yNtf63MES
o6/yY7SXjph5z+2KJZvYfzYGCSbGhsIDq3AXbLj5RpQMF0G5j2Kldwyzlcuv5NRufmiqVa2ol6PU
epaXSO/PdaXdt9Vp6G0YpROTioF2zksAfgh2cToDL6xtFU8ttwmfbybY+9wGh2up/VUQCquYys/2
96kEPzQzxKYt1ERNuor6hS+7OKshY7dqt7FDitzeJ5cHd7N09y6lFDtaf4QIO5lROaC0+z7SbYXf
OzkuKPQA9wS/u0hUXXitNAcnGKTcY7PTU+yeuE/Y9YhNPOaVTfkzi3r1aDZEPcBlpfPE6ISD3XDj
3gWqZ3a2W82RbNqhilHHH85LoCKtGgTNDitURDNs5OoTq8FlghLHQA1CvdnmSCW8U0TQOZb8N+iJ
grnFTP0kCgLURFUxN0N7xA1a6bebhccziFwxDZyJ6JR1U4k251GgHA4cKL146TH0IgtMiP/14YQ+
0cP6kepMkshyrFWjvVMXzzegRrazrjP5os7+8uk9w+K5qcJO7uzP9i15/M5Yp/4HcP7eeIJkgxUV
BKVONp1DZKRAF1g9NJQzu3LJZySAjjVeYLlOJ+iVA6UvhTx9CQ/dTtpLRANXYqKCtnkb3p0r/W5l
aQiEcCIib9pG5VmDbUkSMPRWDGWFhgDqxDbEBgjCbPSJrG51nz4TncBzre2s93dUK/xx3c2V3nx5
c4wZO6qx11EBUld4xuCGYDZh4pUwej8Nfg7fenJe+m+P1lP5c2fIeY4SMCJXFcdfBa9g9OvXAg04
JluN95yBm0YlrDctjW41IqDs4jtigufzwgNbZCnClBu1KYTvvL0/mC8S1RY7L+xM9wv533waRrKu
KMeOaSzZ3ukmASjL2gxwKoX5ZHBjB4GbyRXsC3PngTLqRYG4FQUYrfsTFJzIcEMXNs2DXikPP4d7
R8M3lsCnEMqjTPiaW1OJitGeOqOEtF4VbrrFuc7aAJDSzcaua3zMou+d3tYl1ZQ2BTuM5x66/AFc
WWovq1vhEcUdslYflycoRqqv7WcPl1Cl4m35Yw8KKo8wNkbibnLB0jUAkBCQ6z+dVgKjMOPmSuzB
Lo+nOPTE8/BYYBhpg+bKp9MXpYYLcytItiI7kR7v6pZU+lQTUpHnoXFfd1tSXh9QlFU7OsRuz+mj
2tWAx0+LgegChfBl9TC74wMPUl/QpBBzBitfdOsUe55kZiw/SgqCANiM0mwO38bkOkW4wwMVMo90
y13mQqL1sShlcLi37lr4dOMyt8vwdLPR+l0QKIjngMYFvHPo8rT0nOFFWeAGtEuY2KPPL0d1PTXz
8p82SWQvBxCmvwEx4NSY/70BdSpisk/hD5e/2LNVJE1GJ/s/u+JBlgSJ+y02ofO3QRJZ55hbJttO
ag0otC5Uz0uf6QXG9WvnGt3AMdK1rtWfHr1XO3Ve77n/5YQYsUb4zHssg+F+dWRE73pnALVqq47z
Ce7bD47dti9z96WpRDaQvwuJeATB7VP4OZWy7vOlnaX2GHjTj7Bh8F60D13VcBb/VpDS8faLr239
NoguNa1TTejrC8N7sFl0dTw741gXB76+zqp9U7hWVz/XS8AGhSMsd/K79jbICfMMpRIwG/5TKx3H
ga8HZqdzeHvZWKDEST3n+6Ystv2r0TXUDYuqDxEn+F3PzzdCjSWQnukOW08HxuxQxKmCUYvs21tw
UqrfR2cdZ1Oukp8JCJYpYcdug+tCxCj4/rUIEAKUHnJV5U5Vo+x8Z5fqTkmwsP1S56ori5a1qjkC
zWZ2hzP65z7hSIOpgAG1hcWgdiRwKWnS+QyU1kV9qb6EmIgGF1xoZehfEMCtv3MXQAzWL12Tdxfm
HpO9zjrZqb1oQ34DGC2I+MfcorZFZ39FFX5dmcl9rZ6Ay8f6n0/KiXyFUI+paBRWSS7LEjWJiWNI
n/HWem3WFzrLrFPUeg5w4BP/YR1A0UrAFkVsPdLXcFSJXKgn44cXwVBclhmBASqYs5chsAM4ofNY
Cyxa1OzKAZA44oOX15se3BPGQrnW9GbEOLuoaElpxNSaNVpnFirwPL0znVINjuvt9BwiAP3vgTZp
/NLC7FMg/OMAJdbhY8xs+kojUjDjWNi3502jFVQ8+WPUliicLuyll9KNGWKOzA2P347RzaounECh
GZfLzOnQZNqAc/35l10BfbLLPhfkHAXF9BQQGjqF8PjkJzIUd+CF4UH1qG/zGP0wzoMdSgJd4BUu
DO9iQTUWHROxbtWNJZfYhZTqWdjpjDno2PtjkSuGXZr0RrdhlChpF1YP8ZUKYWOefNHb+r8M9JVK
3RnTWzdL+TwlIxwd5P6hTVicdGIOz5n+ftvwrbW+zzhwsJuAxI/NBDEWCsFVDzOQtsAHExPaDJZC
NL+Dj8Pt3W4tO/W8J15fLYMfeUWL8NENDZ5MaSgIkzaOruVfy6/Bv7YXF5kT6L1+Ld10ZrtB/KTP
0s+ue5fwyRXd8UJHVKutANgZ4paxjcCzxtXFM5gM9g6k8w4PSphx1ESomcEz893a0eJ2PCiZhoqP
RpRmIzXKqMCOtSQq7qGp6LLKB691sE/djJgrfGo9ROFKhTs6WxgoFyCPD1YKMn5vX3kzUPjn77Eb
GUEs1RvaihSOmx2c35s3nZ6mhGlaAtkvRG++UhihioICV0C/Hu3n8sH7bfrAF/PX9Y2D+2Vd6NAQ
AIEPE5r3ycJOq1gbXox5LrgPNrddB0M43npBGHSLbdaXFkbDnkT4GWH+zd0NgDRZEmSkaNiVxTa7
6RaNy24Y3quBbhq2gO9mI4JLmW1GuY9A+aQ2MbXT8hdX40/pOIeJHRvnwMbzYqzMutJ+ObTZPIK9
U5k1G8pLc9vm19VsS90UMZpjU7X8VJfwx9idIyu+YnlcSwFq7iDx94A4IhR6iIk6ddKVkVW5+CMP
k/Y0csIXYofuUni80XzgTIxJbVXnyB5GM/BlOQ9PtLbxLn5Q9VgiA1/B9iD+fFElqRBt33l+bCpZ
VnOmfY4TyMUOzmoZpVpkoQfLpj/Eec5Vyr9OBRW+PXn05r6AttcgmROx4ivzggkrLhsJDQLc15i1
2uDKOvqtClimpaTOI4EcRvnLKxNW890nFZJczs6lWLuzxV6S1UhdcGUO01SigPiOcuxgWg9GmCa+
Tt1VPQAPOsx4p/l7ajE39GcJnUz5V8e17iBgIYNGad+JTZ5zM3lsxuxAghfhhxHyJlKFy/y2g6Ox
CJTT9sByZy0g8kk7drtXT7ip68ODB20/VVlt1ex4PFHJ3uojnIGzPhFG9XX9UuTT4Tta98utlGn2
H7eQItwFM3L0GB/5cDplVWCF177mHeysyhcies8OPfWISeEhXYczprn/NbjAybWbt3V1SkNE/7B8
zM+Ez4VBPLAZmYUq1yLwO3lXpl6DwZLVkaMpZCrRqKvZUxczXsghRVd+EYLtGgRv2djZcnO4XiSi
xCDNkZgbyH8mGrZnc5Pzdw7hb9Pr/c//5A6WcRQdYiNfnuofYF7eP6nZcFpZ/8ncb2g+kD0Gls9H
xIZZS1XBUKZrREeMESVeZ6gZVrXakYyKQi1V2GVGQjseP8DBHbW1ohsHjUEWvDm39NvRLdZqPMfy
Oetj/9L9CwYKqgVUVKmHJvlUPZcCeF7k59poCEAPiMxtfMNOeakjferg5IlvYN1p7TexyrM5rG3D
A6LaIsv3LikLCEyiSpj65sT3eUDswlkLn5cC7YmYBkqXUw5vx5j94SX9Z2EhAXcDSF2NjDgNfECX
RgvpsY71xqn0PmwYh7kGDhNrMCllL1YxDGF1MhDX2AqPqZ1DiRedrz49fjCPTdtsG5v3MdeYjIME
IYMFDM0xQ0xpGOyvQVeV8LGGzeQCqbDei0MIxit0hA1oA5/ofVk2LoWE5P1dxEhYVjRHPJqXCftl
4dJLcZtchuIVjHyglP2obTjeUUGS4RcsKCO4A+ZR7//FTlljI9omGPxBaKqYLT1Rp5bYxxTOcj70
70GObqwnzUyAi4ZeCYIukl6NHrKbdflsOSXY0q3FJIT/KXkIHx+qQQ3gZOBcbwoLrTivRDafcaD0
vWqjXCZJRrzZynQkhMcvS/tOykO7GSiZsHDcfb6xctuPTCMtntm6TZjhB1IauXC7UBJLyRytfVFv
seZfYNsefRnfggFryHBc6O7Mg5tiNDKVcgovUK7OyCYl5daqRCoDPRrWBtwXiyJpzIna9bSst6TV
rTo3YNFLemv2CxwvqU7q0CcJ67qZtVfr4bir+ZNKSzXONIiEkqTmkFbc2dSLcgcusjJs3JBdYSS2
EnFOoxnqLecpVTYgmzoHRfJDCsNSYrPbF0zipTHh4riSNyB2AUFctQevIdJfElxjPQx3XzHr+xn9
AajZ+hkWBV7UgL23m7PqTYE9dTDfHIUHrWuB9kh1xWZ/bDpNBk2OBrvn+4D1/UmyynYcPHnrnlE4
kkawd+D7pzxahXXNwuOIc6pOs2sIpLs3TdQvKDPTe2FKzs1Ro6877sBYGQkiL3RlcDyRMgch89em
mxxjbO6GeHiXnrcsGFCEvDcCnBtP0QN53COYOVk/LXMgl+G/BKVT1CMT9K7djbfFQCNuZXhOJ+ix
plUkHIIWfHW2bU2EUAumOLsaBJ10mgQTHoGR+FbBEVfT8BqhghwKjS23GqjpnwqIThYznQdw59fo
tiezeRRCGjuF/NegLXX6KL9jM1Q1bBt2ATUhyiROzcveS/bt1yWy+HcQiwbNYrUlneRWOSwIgzA0
FXw/W/WzkBIwXAV59ZEitxb4L1PDhE3ZB7TTT0on/9bmM/MAQ9lvQLDEzyrxFGi9xWujhxsIQHC/
Y6Zb8wzMFHO96xz3t3VgqwGg0DLr0JTllnysNkHSXJIfWIVshtL71WRHmfy0J7IOjr/Sm5MnLuFx
4mjrcmIEVE5CTHJjjZWf+Or7J3c6SOlJMazwG1/KQ2l3B+RY2zJ0uL6fWjr3W/Eg2SL8J4CFbXqI
vyn5CH0h9tkmG3HjRI6S5wQhCuPMlvwflB5k44OjMVnvZUgSer9bFyzmUiVrGwr/XAV1ye8pKIof
KGx0kYeEz7vEwfR7Y64Q55MG0PFkD+pXAfBYlTK4vGLEoY7JLOHm/kvBOQkHZYPEhMIQZOzSe+K8
I97TQgIc2Kef+moKxTjfWLXTk5bQij2g2z8MWcjXI3VU7GV+mmzp5iIBkMaO/Klz0nyd++FaogrV
FYA9sTyw6B1ZK5w6KN3KNVq1lcrVj14KZ1ajlwQ/P/MKNrAeXeINyxX9adM9PX7Kj1EYFWdnkDX0
AGNVEBxndtSCktxeD3UGV2PdUzaMihVnZ8jvlHCQtv920n5cTQIvdPIy3/L+Ip+xwxC2IiGoKbYz
8LZx6WdBrraQ2iUO61TuMmkyH8gq2vYVWc8cSir6GoEEdMnNIgL6TMJSvtfjzRz/SkBBgeYrcf+x
Uh5M5n9jMaT/pa3mnsMeUyICxuuXUplBBASQa0AWTauptOn07ZDbNVTQwnSUN+b3f/xlfQ6YKQ1w
HrAj6M+YvXy0uwmIIs1xSAeeztxeNP7lStvQ/fixOjoBFr+SrUyIm4U1JR3LFIikm3xITE1ZQGWg
Y1BKkdCeLWYT0jSCH7b+tGbf9WHKGA/u05KOuIbTr4BTDtDCS8dWJu7PEOnrb7bM6t+ZsHkfDd1l
oB0rGfFmIQ7GMbFKl/SF5n4YDt31JD5gmTgwLFhazuhVaFIS4yD0esnQH4YP2mFxQlGZeSdKxiK4
tnOeK4s2IMRl7ZDdeX4EXnR2yoQGEgujg+C1lgeWK4uNQjPsKvhlp7tI/EDV3C3wdenubzrF4IYt
4QCnonDH5CKwfe+2ROnNBxLMuNrjU1VMLHyUDrYLexCyONgw7bls3xjxCp+l05p0c/ODCGpxgSWV
85A4UpUwozM/8gQ7NOBXa04d6n6UyZw+phrTECXJ2ojwxnKiJ4rTLTn3A/lvoCvutwDE/MhVIr3s
rbkQjgY8LILJucdOgRTHbKBCcDajP99T03mBzpa6I2oruvttV3OzhZnDG/kZSKAnHWVwN1fl6Vgh
OpcGfB5KVofTYGltydoLjaL1kfNHlrbjVNoUo1H6Q6hYOL2aNl1putSYJcsAn3VDUE2lrMMbN7yY
nzZcXD+jyaTrQDOFFM1raSyzohjI9VI3VfKCv3Xw103MDJZ4HwbVimPL5PJVE6Yfo6C169GuU0RR
AFuNdQfrys0TwIaDE1YF6Kr8ChWDlcOVN/bZFvsZh2VpYvIITSgJBfBkxm4/L45nRUhaLVEsOSC/
vLXLwF/H/B/ZkCn1iBJ2uHXx6aBANb71p1HWQmLfPHmUZjuqUlsvMGi6M8XU39KN4JtMWgWN+wWm
vWbKhE/tC7FqwF2rOGnzWrix29AW5rTLj20FS2Nhse2y05uVm3/+LnmFGXa1CNjrbCcQ3xuEhp3S
0FSzXRnWAvg4FTbUm54IcCNgUTDu5g6Q2qAkd8cYSucvaChwf8qoeeGLNx64+zqb5/eF0CAVNGQD
0bndDfvZvO0nWN+zccPyaU2qX0kngdX/6DfdYjIkClMzyxB5FmKcxOVaxdZFiI58He5xJn971KRO
n7ep5UwgEnhmugU6g1IBudjYR1TgMqGNuhsdWdEtncGak06a29afPZ435deoDtKYDBzC3rm5umOx
QjrA3i/0HNrwk2gUojagLI/+1IwyFrxzU50zM6Y8S0nvj/9R/5BSJB2S/C0sw6UCR59Ev//Cfh+H
GyuMpjqURM+oggG75DUvaqVw+8ThyVnM+rcdH60ShqJJQUtXfKc1bkwSFJjFaRDqOEnsmtMzlM3c
+ncjEVfSPJ56vDeVbWjXfLRCRxSka+Go/8iG4FEjPEtzA8gObMWaeTtbzyJPfHK6zzWWsE6hoGKW
KQRIbg0xDHLd+8fs/L1UNM/OfnIO/reYWSZfCY0vmoSFwb5o/qAiAoGVgYFKQtotABWViGWM48jE
MCjHP3LQU/kAvnb+4/qBwSZICS+M/SOIq4VqAsaG/aUTeZvt0d6XCFuuG7TIBHNHnh0RGqwffd8G
gsPVvzYPc1Vba6g1/niNJMQkqDy3IiInC4n6IGVdP6gS7IKWGcweuXKC1OV++32BGJcn7fD4EyUO
SiTYGu12X90hLGjtTLLyPaL5mNkr723nKZyAIovLbsUaX7+o9xeo/GwmcSSB6PW38i+lvCWuuTOC
qQtNdqGeWfg0rNHB0LANnOaLU0j+Dyb6FgJ53+BTMsG+Cx1lzgpYcgJ8KMGy8dtlu01TH2LrSgtC
DrqWRg58HVWJYIGNev5D3CPMoY3tIXKnvPFomfYZpxp9T6/IkZxnj7BbE9CuuJCmcEcP17k3USu8
bOGJcvmPdjEN3E+y3pXYIPb3SOODoZ1l/f+0uoIjywhIsLg/wBAv21ysj/3dtldyw1J+GXqImuRH
Ek0f4zjs5C+o6IiRwwXkQxatRMOMrYGRdV/GqH0z7h3AS6m8jU/uY/v/Oveuz2TPTbShXqcFXnsb
VdREL2lHBae0elZclqdk2ZgHKHbMjsA7nyoNLYBiZ31iceZleuWMDF9gSgled16ph6kmbiEhJBvp
93tcfLf3o/ddb/2a/H6ZprDO36+cJ3IgMQvQFjtR6QUXhz1+rGs2k7ZQl1F87RJthtbdywFs0K6s
cBvzd3U3A9oYtHYBcuZgeElyPpe6rvLYg2qZMSu6WeeC32sOsPkVLHpBWWtqJZJx5zfMdg1JbT80
jFD9DDwVKNraBpmGTtGh+j16bY3vfpQSbNFNy32e5o/i910Of1W2orVhnc6+0sNtPPwZHTjlfaF1
6UPEJzf8Mi1uv+gqS/tCha6Fl/r7YiHUrF5mQvt/89PO+ti6jcE4ev4KpXw6aaGajpYVxWTosInB
s12sdJAA2dTMNn0pEHoMjmBRBJQYl9rm5vxKAHfmpCvlX6KAbOrjnPKsgdFVJh5yb9Jk1C9jRAsZ
q/GzUfjskXBIUAHGukv8sVDLqPgvEbnv/Oxn1DcQtY+ccasTTbXdSfV0A+Gjix7n9UsNtP0OMS1Y
CcGLWYrFGFrAE6wkPKZlHnjKHrbkRzvGgTorqeRiiUem0sqXfLDjgf0Trnkz5MBgMfKvTd/P3g29
7haMSGCKfIZO3WCxlRGlu3xLBChHipTKyMNi+dasCCHOBFvHm8WWEhZWQpItVX6h7Q1UCJtplMsv
x8he1TYwBHc/QH7UwjpybCFPOXbg3qjypCQF6Q/CxzfUOGpCeT3aSdFitvRVKrXI1Bmwq8E+vrEQ
Oa/llppa3954QopXFBScb56Rn4G0Cas+hinBrXxXc1DSwcdHu+qJm3ePA1BGFobpeCATFysnbvUS
Z7zHc5+1oQ31N/nDUf9EKHTeJQYhJ3Be9BRyeii4LO9hC8HUaz7C+C6RH2Bsh4znhNvL9k3uYcrv
IItafSXZEkUCfvFuMVIP7rcpwLz3RKALIdoemSbALChHmEkR/hRODOt4oBhljQiQngMuWxhiVHTm
85nR9kBpXXCZyZz07qbCjUIbsZGwJVnBAyXpheNNArnkvdgh4rPBDRvCYoyzFXYeodbUKOg6JfdB
ZBUrn1GkHho3PV/YxMivCrfnMDzvuJsk5nctorieWWeM7Sex3EV+n0RmZlPYATzKLVoeHpF47mhA
ez/M4jiUal8F9yMAk/rpc4+JuviNmpsBQviG5bt6R2J2ofetpvp5NtqnABK7toQ/7RsuzwZWdIqK
UouBDNKvKRuIbP7Cjlqs0u3OVNw7MsB0RRiz1hSClFIeHsyI+rJGFSmxD+eoK7uDlVWK/FLGgvtl
zlQHyxKb1C4Krs/m2u1dpaAm0EncRo3ert0xyKcO1L9n8DH1dhTdylf6i2AplkZewrZ8aiwhnnss
iZ/4Ptf97W6AoYB6QOAcHKbwjciwJbsMbGRkf/I9mlqUfn/qw6TIWkkpODZD+EL1CILqO61y8Upc
uIFWmx2BzFSAQm+jmt2banBRxFMPpBjaY12enGYxxRBOMzXDdlFuARTd1dIfjD81gybN2V1hyaYO
LUiwB7crDJi2qrNH4WyXQ3Ugxgs2jOq/7p2+DZhROPHeFs7iICpR8XSO30jaU4ktJdhbXPjr9GFy
dzdLTx8MdMaB4dJD3XPHa2liXf4Bj+8jrjC3VRuxIKW+zbIy4q74ohV6aP0gNolgtoLKwsUI7ZdI
JvMcQqdRQGbj1kWcxK4ZVB1FDlL4vo1kgz6RDsoNH3Dzx5dzbaDoWa44RcY+1n86BJQkoJVKv8LZ
1qN26Oqy8mb/0ZJvmKIRDSvlsSnBeRO5BXCMkscEPFS5xFwfIxsHvGhPAeomGtyhaoUFdOjOslPo
EmgEe3DzyG8ZkbvhqiK802EV6jlsy58hx8GjKrv77plJ55gKv17BuRxKJBzG9R5K+09NHBsTwrEi
jiLq3wTma9pM4lAtKLxA0YK3IVaZyPXgZYaIpBhphy8L4L5NGf64Vzrpan8+s94EXLGCrcXXB4jt
40GDdyT4Sm6RYSHQrWP2SzxOmnoSHVlFBU3ZPWg2tpW9o5vMZ/m2FeRFMp9VpbRyQ5sDGy3AjIEH
SsXnscpyvEBo17JiiM5kXCyb8xa8agt1xBxMUfJLUVKDo9FtiyQkupLS2oYW9KAxbNKcdfxcWEMA
4TFsKbE32E8ofHuFIz1prI76WqfP8S/vdFww1t1se15nxW8K0vGVSNg6wkQ0WVuKTDjoKvURe8Tc
UtAuPsFBL+OMVlsFzmXfS8hxQQSZGP4angUuf6aUaw+2W0xFm5bt0Um5ybl+o/Y5tfGNlVWsy4kT
KCSLZjG404Oh0NFOM/TBOQaKfqkst7qVVblvL7/Tf1wHFNQc1ZGhJh/mN3dzXLUdWO1sCGd5j2pa
lOi8Z65flW2I2MhYq+KlQXoySzLkhpetbDhfxDRsviPTwRwqh2Fztv3fQgA3ggYOTGW3Vv/oNQpk
ukWxvXc2GN1MLp+AALqLSEe4w552+Wr6W77OZi1e8gJ4747pDIT6qEYJNyPyQKJA4kkkPNIANHsn
Hhis1lg8UFjBp63ZQJAotwuVpNi4qrpVw/wpE3+QSiTypabB5Egwp5pk4wF1UyQtEb0Lhn1zqH9q
gsmOrR5Q2yFdT5dOIieeHk8Gem+0uK7Y+QMiFyu/K+DTOju78eGHNx5RcU6nj0b0RLI3gs28JDvC
hFYZT7wSXFyTOPJF8qWqCT0RlINTmFcrGuTRjTe/+l2FGN5BapYzROC7NB5rNbzJnXSkfZMVpxEC
999q1qAJtj2PZA2kk4Vj2wFWOMCcE7kBWtSQqfMyxZAEdrtqSyDKIzeMErW9GWEenvabbSsdR2tm
6vdoeokM8AxurH26aUl/KWOi/HtmL67RdujVOUPw/5sNCt5tT7KtvBr8lycL8sGfdF3Cng5zUk34
kjLgYVNOgV9fWnZhH/fJHQD7EUreNwRolzTz+NA/eVZawASFhbk8IFvSz8MPqvgUAp1FoFJztjpk
SWj1QC2RDo3+Fu2mccSBr0YvAbpXPG44oHcXmJc7BC1vpVlJIKVrlX7J/gjS1B4IKkxFPDkzj3e1
xxI+zhEDBdnW3t/o1+sQquek1mpYgmKIwolwi3uNEQ/PfF4ck6Akhe1+kcUI2dJSNDtNUKTgn2cY
DFhD1N42VHJ/ipUiCaLL01hvHYvrLX882q3kjK3EoPkJHQ/XHl8BWb6Dhhn3mPjUBcJLpK10+f3y
d7oHvZ6t3E1JorVIF8us88u27vluKjuSSR82BH1qfWRt/iE9kkT9f7zlTC6PQH017cOLedCl9i/z
316hHHEjFdk5rqTV05Fp8r8T973Xbw05h6+0OrlxZF0SEjguOTQn4fQiDJ7dGOu1gA+xtU1h/NpN
eYsxEQSPa9T1jQSIMhHlNj5A26p6hXCP9+AMxKw3cg5+jT7ZPK51A9C5UhAKbSk36LodWMGuozMR
kGE1K2P3PfXLelM+GswwKoJsQA/03lUELT2f5Mxw5wmCQUvMRJrHDGsiFaJ4KU8y5WU3I10gdfO3
VkG2bW/H0e+0mL5kkwDcE7qih3DAHzxBogWoL6Cee0KEL3IhidpjokY8nTA55166ztt9X5frMjLx
y46RhVGIynciaGLnC8R+vvgVZj/K0Wl+E0JbximwMmBrzhWzR8IBPcSnzldCeE6tEaTPZ2+mBXbn
A+pvZKsMHlUb357Tj+1Gg6HmkUezn4mAk83o+xKrlpyP8egCtJim+QfYR+qL9eC5tTuGuzc57YIk
YgJ8k0ESsZ6RZcToeXSH2d1L8onb41pT2nMoVxJbVGlSKxvv0ojdhplHATaVYqXKThOlCOTAwMcf
Vpb76PNhm8qAsE2UtdrJajf+vwBRS8Y8m4cUjWZ/c17nJIJNnt8XAF+HeucFGYRFUfa8IULWW/LA
Et+dmRgeg8IaI+hy5FBtfafAAm7Y9CISllx6jlj9ZXDKkyeODL87dwZsJrmboCNax7xxg7J8o6MF
EUnR8zIu1k785B+5Vu4n2L4dvKkK/TpFfX/bYFTehSbGZYlc3FQvBXSH0+y+Z+UmzbaDU++6/G4/
BYrMg0wemB8dJcS//7x4x9Kp4JcTvAcfx7Yikhi0GajlTrcIdpg0l9Dn1zFCj0KRPY6YIoC0byDS
TCttO0Xed0fb1sf8jwr5h5a/z17oP/f4rM3KlK89WmhT49Q+Zh4f/O1BEMhmwnD/EZHqkE+WHPTM
IcZJ0GYFNBXd9u/MIpiO+v4QswF3NECohRtpW+Xt7aQEX2OWmfnSip5xhLOs0Fv8GdxN2NEAYmTL
4WYyZDfsEgQJoQJfUwv5KIh3wNMcwEfdF+z1zkPC4NstH2ohbxELqCqbX8ifZlGYHf61k+BNRgFO
wAkrPoyTfmrfqziUT43LWm8RNv+MClyyTWvoz3H2Mi114ANkhUuSz+THzS0l5JA5hdSda30IaVtz
3WhZV6Hq5frsk4ABYJ5Rwo9Dg9z1Cf9pX9ib+mvZquA6hWhxm0ogEUDTSBqJoTGQPev90zaeCssE
0f4Nv8DgOH6CvcGvVY8oRw8/jlY9nOxY8UbPCVa4V/RawhLtSKg7XCzJEgEKsAyPgnnn3CY+a5LN
vkedRcmk89SC9kjgwwwU5pZObhgoNNgPP2Bv+gIBlAZ+g9rbjqYKnto874Juu6T9fUtDURXebfsb
xnIWHkFkrdTWa74Rztyz3Kt6ewYDS9J7VJwLA6JyC8hXAdezVUwIgglNsIlSDKziqSXjGtfaCViH
NOJS0zUa9SVzfjKTBd37+opMgu6Urp0ij6CJynG2Ot+gkSyoDyWZstOxcqeViTt8fpdUUxz/s/V7
MWqpl3rUuJRjKp8vG0IL8z8cc/DnOoMPC4O0xA+mMX59stELy4NBcbZq25GhGfvjfREhhYUGNtfK
uXShEG8hm8nZL7jAz2kplvyU0bcMh7yGglYdkoMcy/dXvwr265Tcx1HR4FfgL2vxs6HcmXiV3RVT
Av4fUh0kkgNvj7YKTPxVH1yzRDWxF3WHJ9C9QBrjyErHoqwHUImEl8sB55obaIc0GDTufkxTZUm/
MsqX1QxC8zdz5RNzzl1TF3j5VfxcQifXrADBdmhhOFz4irO62u5hzcterrmNTheftTsCWEHCgKht
ioZqwZejfPBXcNuHqMXRP/i4aLqKy2RZ3zzvP3sdzYkeO/EzIFZLH6b0j4ZxJN8AxGjvgsUTK1FU
SQdoTz0SileQH60j10+PKj5slCN9iGOy961BBJs6jNQWn8rj7uDePhzSy2HeWfmY/98qI3BPqdRU
v84rOIHQiBXjnN/A0XEftLvGBbsGYrwTcKLHSNNwnvLiaWgVGC27t2+2AIWzjdT3mWTsVv87Xv6Y
nyNE0Zo9Qh2nHZcBemtIWAm1gH8DFDE9q8C7eop7ii1uOVxatyXh09gXJfkCYruPf/Ur/ixazBZV
uOPaghJiwzheRtFCqSzf6M+lxHgfQ0Xs8WU2X6dZ8SXyvFN/mUsFd++sX9D90P+K1BDXFZiBysq+
U/N0NJgqTEXsklhOr056EFDFgaeNTExTrkzVQobW1pgFsCrHAtAk5RgezSWh8BCF5ieGQkWVRNIK
ujC8/8cb9A5Mqqzph+/0H7jl36etfoLu072tIxwvvIO0fijB0eJYTRu9r/tlQ3ZodFOLTmKWM9Yu
8YhmCcs70xo6vzoYzHFoQMrt8YWn5dcNwQA8Q2dG8b/Eccn7lG8F+yzxD1OOImct+0dQVi5HrjXj
7FK+BlH/XtDIAuL3l34CtpRdJN4FcYaLi7fDrZ/PUeFI3ESsHgyHu14IMU2jTGGULxwTMk3CpocF
bOlMfdN6m72Z7vY2BLLSZMVAhZveBzLmViFi9rQKdS0Sg952fGN7VjRLeWqNQyx6SNi+XqisDJgq
iyVDSK8qIzyI+t3sQqSMKkDCixHi96qo6/aszPKooqer5rZ+FgTAG/j2gMBpz0LrMa9aY+S2lGbV
PZ9+b8MEBMh0gQe2HsgFXgcmfQQWdjJmcHSKfce+9L3T8u2+jO2gay/a0dPiyGm/K6N+J5NnhXE0
BjpCDjzPM4RnKVzRiAJb2SF3hHGAWcu5E1b53848O9Ms2EkUruAU1Hz8b4XoGDE6E6TZQ+18dzm2
gOZRMAd1ybpIXWrKCPCYnlHmQ34LCA0EpsRWnxsC4cNVLlIxkV75zC/+SYABBDFKzC4R5/hP+s16
vLy3UrACMl2XLAbdVg7mNUCcE2br8QJnuykvDx9cLk5UhW+DRN5PO9j6UKyh5AWyNrMMBjTxtZZO
u9SVkkDbDpgdFdzQSQtWAwFOcLCDPcHh6I5nuJGpwe21hooNIXMtvi0g2+EpO/u1Ct9rRc1xIxPr
W3c+UnbIIVNaJDVFJGcI1VcbgdKwfsCKZuf+9QTjt5vujDgtSwlJYrnxVh+urIvzQoYfnm4R36iP
S/RbEOgL/RvcXDt0t1NY3PrefU6faM4G8sXzgjSh2ijN9Xpnt2II/5YMWrHxs2Fjdu/MFsa1+yFA
KggUE8naf4vm/8/M6p6sYvXpgGWzaJpE5DC5hzCh29h6Ab1si8JEW75LJYVK+ByX9iips7K1hKO7
OZsC9nn3XpaS4ifM9JZa0p+pTgp2RoJCHbdrXxqoBQ3juaRB+RzdvliD0LJlLhKv9zHawAeoN78/
s/WL9elBQi5FQAntNDKJpdLZCwPgAK9ruIQ3hWLGY7jzG9dwPqPgTBo1CRo5f46Afn47jc/KHKdO
+SHglyeDBd0O+xEMd0+X2HcZ4ZkWGmt3R3pzOVuC37OLlVH604+jurXgkdis/NHvKNMbZECl4D+h
yFusSq39dULu9jYyOP+Fo+VMsGGBOj+6xQk7sZ/muqI8M8rpJRAawLE2X8VyiIYB+vcoLyjfK5Ue
t+di+i7XoRwXS577+eyLTBMJg+w+x4UvC6NuX7nxL7SAVPNPNlFlRklh4YcOsNot5fI+YE4NBFKT
eCPt+4QRZSxpQFSpjRdmmNWT19lAzfOjXwURyRm2kz1ZLu4hL+QxuWXPBPGelT97WlQ0XefXzc3L
HrSJLMqG2Q63fSw6YNZDXkvXdSZoPz+WVOhDc9ynXJcucobjDRCyNWODTPaix1bzHM65CQii23xk
J5kKQ7hWnL2QIJgCFN/P3EGhAmqmVJDTURhnv4snQb6SlrlQcGIR11ubr1BiMuhri7lkPsgWIZyL
RTERDVOVD1SCWFhypW98+ww5Vbhgd7K2LKZqVwaavrG2cnCwgV6pTqmVd51Xgueqt53uSjKa6vEa
hWxJ4DrBMrD/Z3J77W1MrMlkwmV6daZ1NHFg8nfIgxvpL+mbgIn2iqsBRrEGaQVCnzrsEgmZqjeO
nUJlkQBQ2FOweQzb24dAhkAiEqhQFMXF6XUk3v4fiRU2Mk3IKgdwOEZ7vFGFhgKfo7APC4lvXiV7
XMa77Oz99fOnxn5DQcst7X7+yKA0E5gmtu3aZxMLq2QZpRp6hUesWigKz0bMickiG2sOCoXpRl1d
bGtWVUIKwc84uj0g33A/UKgu42DrUQalKKDXSx32o0JsFf0IKBok8im8DZoWpYH1h5q0yjuJxeLl
Xkco66O9dRlQBmxpcVMcN7HCFxOOdqmHR713rRKdtbVDLvO417tgN2tJ5VoB/WeXmtWTsWUJpTum
x7aV4wyp0BVNbkpE0+hV5IA7asmw4+RFcHC5zjHt4Xd4gh4IbtbO+1AOVMgma8vIk9+HgrrCmE/h
E1DGA5PTKimcVd7GO8nxg/qmPp+BtOsQFWSWcdTw6M6uLw3SxO0duZ3RnFh8gIund8ddoN5em/cz
FDSl9oqi/YvuEhYV+7ds2svyJp4Q5Yv0RLkg5VxxvU4RKuv/poDTVPwAbmke4MFosQZ9C7aS4i0b
e0o1evJLt8A/o12e+b4mSElZnWE2APLY9b+lgR50mp9cvTTfNARtYeu3YAZ//mNGWv/X7ug6qhdw
oFRH61tld9pbBYOHuxCX06UqnpUWgQ2XedSAn9I+kDsAlOip+cZeDL+gKm9Sa2rzIJ60iGP+3kek
stJr2U1JwuIpzq2u1MYAfqP2TBdayCDiZt2LUYIDbVODhNWts7MeHwXSMwMaFpSCylX+ACunbkTE
74RTyeHgFDvC9jiLLzKRjlDPzISNdMV2Y+ULH2bgznTiUFlaaNW9IzFKWYFmvbYoQUqAU2NnaBTY
Pk8yq19yTkZcTt0YtXnC7y6en/2NfIKd5FeIgbclqHcPVA9eHbiki+PbxF8FhqX6kAPMPLwb04dI
MqIiM3VOFbfi72xS/aeTrreinC4mvKzS6ACyqEXsq4eQ1J++Melc+U93y96+yYeViCSzOD/oIiw/
3pBT5MgeZw2gvVw1rAN43TxOfqPTB1iR8+H+GHs5toFFJNPyij3S7Hf4vcHV2/nsnV/Qx9IcI2HL
DMYqN5g/Ql4glS+qq8QS/m8KlfUimyBpLfcqAR78FfosJPLyXz6v6AgNn/96kDha16HStRBPOXRI
rJmwhenkVjEbukqOzTflVCa+eMKdnVqLybcuozXHiGaW4M24kLt1x4lFIOPVd/jXRuaVAiTKNPnM
b00UlDhgcdAqJ2CBdLhhDt4zESE0X+1nDTjjJTGXq70+rPJ6tpDtpS8gI1sAWYarR9Cb9RML5wVo
cZLrqWo2u2xQd7xgtLBUQ5+T6jAcBS1obsL2rYpTfXoqZhcxIdpA05gfkRSMwZgPfvlJEyupUowh
YeRCOHclcVMq9yNY0wSYsiAtuxidvyytkVi34A8kScW0O8zxs7+hK+Joz4nJ+seeeuz6A/LhgCaT
xaVPEyX+WErrgLHoK6axDeXE12UQ1wtlot0Bh8ZqI7n6/kOgbDnDaY3z18a+QCDgpTK4YiBToE3N
NCPPghpJ+xt2/iac+I9S9kZ03Oj6XNXJV8mk1oEVvLuhiHZDgs68Rs26+6F43sROVH4Zo/kpuWy0
cb0/8q0Ydk4RD2AewR22JRzQsX03O3IjL3l51wgN/ojSCDiGJMnKzAnVaqZGZiCvv2+nwmzG9q39
ZHIXLR/+ZAjmdKTVRFm6AVbVn+duepMPHYrU4iEDU0Z1diHpIQXILPKvJlslWy+C4pI7qEgXcX7q
EylCWHKUy+WxH0cNl7WVOwcBK9/yBtVKvGL3eHRjZls0tGnlh5OZee3OezE/oot95em1udv3ew3v
RUIHBEh8z/0F2XW+YlqWQeBMYiYVmGqdH3ZCsBtXWP26KFXzujbHlJ+RT2CZ1ptJstr1Q3d7EfD+
Nq94YMWdLRkviIiqueV5Ymw8auRPOkgq5uatgqH4UWv2vNzo3su81IFjxhA9CZ5450cxTW+nRinL
5W+9F3XBPtk3wQrDsrojSC41+GGbGsz+pfl5XUPHd5JJc+EYYLBWbMcKILGQQ5VJIg+NfHPXdhZc
J4mokNXNAmC33eXv26Q80SoWkBRERUXO8t9cD25wJJT0gFWdu1N6I0rcZCgxfhT0K6UahnUjVhwY
2Kx08v6xLJ9TXqS3cTZlKLm0DJ5NX6MMUONUSrEGHaD6no/vtEdyWSTWP9MVKfGqwwxmdPb/CkrT
zICdoXZk0iNJLzSGFnf6P5iAFe6ArtA99CfjxhqMyd3z7BrJYrp0hmUXU/sIu4qowCjd+RtQ55bH
V5HaI5UwaN4U6ucFZembYspk5Dx1cgP67FSRhZmFVjVcOd40n6RCRBpMubgsaLZ7NER/F8geGsX6
N0hmtnsaUCdX4eIorLakUgFmRSJXNm2eR1dOo6D7/mwISrr1g/QQGXldLpGp2Rbu594PMyEft9mE
ILgQufvnebKBQyA5pV+mn8gybI8UdKz1qf3pqXk0vu2Ac2Wr+xjSP/DXjLAerlbP7IOZGcBPtvVX
UZUXmnPb3tKuIdPxBXGQBFVyw+UdMEWBir19QNnxPgLI/xW1PGmy7WYnkEiEQtE6bNQ+II3JonBv
8EKY3MzR+KI9VBxmILURmvKDtieDCSN6D8E2ZCi15Jj6NfxXWUU57NP9VTaCAFyMPrpWX6w+ccXH
dBPGuwuXQsjTpdc/ZPRkDy5viwu3SOA6x2Vt6OJIGROAM5YjTzu8rlXS1Mxj+RkG8Faj++HimQuK
m6FMLMKXKx6+tDTrZz/WqB0D64ppsjRhD0cc7Izs4X9etzjDF2kxRRvb2ZTeW6rcZno+R/AvKwfK
r/YrqV7WvuJfVs2NnuuGppZkW2Ow7p+QztCbERLVSCIYogK2ZosPX8/+kb7E2W7vsmeeo+CJfA8H
XiAC6VSIyYIdK6e9+c6Cn5zumV3e96YsQ73Ul+3PdPShedr5Ht3l3A3Ykzw/RX1OsKzl2ixyWo2P
cEXeCX8+uwhW8dUCqbzONkFjp1e7jQhqCMqbHFly2vsGnZZ7aYVlNUq7GuaxVS0DbuEH8XTHAmZR
cn3dpUsGAjM+mQogUHbM+SxPX4xLdUOt3ePqk0FNRUGfY/JKYXHBfhqLFE8PLmGTZmZjeT1vHmT8
K41vUibeQ+1USmDa2eOUyGIFeSz/otPZgBm2QXVJXOJZKXaFu0YSGAl6Juuy+qV7ytQDt4uV2aDX
TIb6mkONYmrOQrwDcG6AKJdzmhfRmXfqajIWYutceHNL5gzHHhoJra7xGQeqG6cbG8802RxthtiQ
emk/84MsRPwYEC6RFM4GEkFXzQYcrvX6nfr1HIYrgLZ67bQ7isiX+TlzmgBr1AiCl6i3HjSMJ8tu
nO1RS1QPMfNaA9JvTHz8Az4SAcbnBpOZPdNq4b1UpqLXVXgxQcLL8RxUijpAIzypj6o2TGSkvUqf
MMLCzkaO63i+aPlflZxua7G3Yx3q+OFm2CXxmTBdau429tvHlgnHCNTa+hcuPw0ZESkwYK+8cYvN
aC4ddFf2lhg+kxRB7NkBbWcI3kqIdYX0lZkf1SikYtIfg6/CA7uQtLtXYbE2PGxbTIK6rgXSQL5v
Gf1M/iRrb9V/4ygLpivX5KOBLHKNGyGIQTyOK8XSVrvl1wgCMgqx1SmgPLtUieC0pBEElzR25nor
OwtW35X3HCjTKj4cObxA/kugrVEOJLGVZsrDFez4c8Pu7uhFLpal24ZzkbEALJhXxuD990FWCq4L
Ab+bxi7rrEIXlX2shpUeXPadsr/a6J7P4mHU1vloflwO/oj/q+m/YvooGzp338FXn8SIVJXrVZyK
6K0skTxPuwONGndzZdYxY9YKvqAkFOkVPIw6ymQMVEkHta9AFXKTTvJWYMaT3mQapN1P43UApvFO
AUemKOYBDFYFheQrQeMAX7MoUZvyUrCQoMpmXohUaXAjcjgmxZYDCb5OqpT74NNH0IZ3cyBuK0S1
YkIaifJ7qORi85SrAOkRIyFNZc07zZzv6YBfghtvVjvl2blHmRWCyb1FxvJiFEng9volugB7FhEW
ukfj2bB7xmlJfnhtYfxsnbnyjMKTL6nGoAHMl8Se5D6xawHsb2G4yaN5wcPTLi8l5Rwgr/STk5jH
mJG5WBDNE4vv8pECkBXgnYCQBunOhNpI/fnoAxh3g1F0smi4dl4Tou+P4uYgIuXVAs2KOI4S2BzK
yC6JGewQEIMaXPDkKMDB/q6tJnzChC04X99feTGL+kfnmMz/OX38fGstCAFFfpqOpkyoc9xO19NA
FZoZTDdNiBojAiGkBUsZSqBx7O0RiFrr4RbRcIsftTElLWgeKaL5IGPIUnuMmkCwPEJjCWgnPmer
OM/xcJrOZKvXyDto+f4f+QExKIN9ZPWMbPvPoXIw6csDl4Eps95og2RwAbFru9uvsD9HW9zi9nzP
e37y+reOj2dP8C4U4BZYehTdIvHLeGr0Ai+JfjN+xbdei1PetCW4EuNsCvWOPiflCXF74FGup9AG
LkiJWRVxUEpNMtIuD7Y78o3ed+WdhoXxbePL5pV3vVlA+EieYA1Y2m6InaEvlrXnluWWKq+TDAqx
GrQRhYpiGlhJMcueLi92ESXXN/sOEnIg2lACN1dA26fzbaq9+woNT7KlFeQog66GJRSg/jXBmsAN
qAp459RQ534hd86PCLVfvkkUYFj2VfAwbM7hKO5JZmOWgkoaVxxeCzZpCeZihbTCEMOciXVpY++y
5KF3vyHhdlL9bOt8TDOdGAeFm6z4vVmowA03+I4ipKONUl3byNyA6eBnwrziu61iDIcLR0lBb8I2
wvZnSG4MibhJjpC1BCfcY18T90e5R90LqOhPtAFqUPmAwqjvf4Hrd3Z1P594kD0h5rbBoYeLM63q
VTsiaGhBdszLvBVsiMLfqZj+jzk9EZVMwtvCtJOBF9sOSZEMVK9lQvp9L+ke1IyszdV3N1q6WKUW
qinS0HGccGnvwBDo3K9j+AyEAZiaq/1QeauAYflVWU0u3ZY6W0DfSMfB5Ro2PtuCsAJYWmnB2u3Y
TCcqnsgENNdG7BO1iXNt8r1dfh4eOS57nl4h1V6/gTcacv7q9i8i6m6vYvhfbDRsI6nM78ByY4j9
i5todZtRwxplJTLzRVizLo1zqxIfWmxMKclGyoWRxy0KuWKTatC0azcd8Y4xQQ/nDC47zYCttsN5
AQyllyUlXlWALADsn/0eoCXz++egD0nExXVZ49KLSTgsZKV8wYWPJ6DqiWNADIqw18+yC+T7MI1w
KF9kfY6CbR/yQz4l3KE2l/syKkoAalKPwsScGD+RTpp1hN69rD8ETYxhNK7N/QMbbqBIekSdKjlk
rXLKs23U/EjHLVkBtr/jbPj+3nPIEaM8bES2C3NzpA5w8DFM6wrfu/QLyxdvXNw5boFuEn/R9FAv
hJ3HYGeaK+gSTG+uunMKvTzk3zC1hECdiIgOJvo6phVDf8ko3Ijsh63s8tghb8mjLrIyDTLQzbX3
MQIjYBJ3dEs5IiIbOjrrl2QrDAIpvsKoG1EqmZYViNxWPJSPFaA7UxzwMucT9hbqO302IxChmGyg
ZGFHQfDxGdB5QefpBF7jgREnqJg6wE3UqUt2ss5VFVjw2sf7IdJXFI60XE89o+8QVJtgUpqXErXR
kwSm0Cj2H9Yudnf+ivr/IpDNW1MDc3Vnwe9PC5iqRSPbXLmkQCmJyTz0zzy45vHbcY49io4MmVwf
118GuOKth9K68+BSfXRE+WB46xuMWqcPA9e9BXHczgBJXVFtAeEqcHFIWOkUgKN7iASwcdJ1b6hZ
LOMfTcVXIIe5dDtkPMpKISVGQnPq5JkIXjkao2delndk9FQsEcRbnrOd/twWD/zkzhujP1C82tca
xeyF19kBvRwZWcwYb49g2KOEiGewdvCW6JoyoceQenoicG69wkuDZQjSuKsxAnr7j01Wtnzi+XJV
RI42cdLSt+MV9lvPOCrXJ6KJ5GTmKKQezcXXEKgilhXCKsqC+xzb/p7xLHsycrJEgBTyEwbmFhAZ
3rgI1SU7bGManMT2Gc2Oyc1EZEE2R5YMCugMdrlTDpkrkrvxB9+jbsf5hVuZZDvgvDaKZaaFz4Hi
Up/fq+WtTWqTVgt2fLQWywnzZMlWyj5vQCeZ0cmlRQQYxjUw9GaqF1j+thSGWe3DuFI43xV8pgS6
uBuxEoWes1Q8BulzDr+ogTtty7dbdfy/LsU6wJXBT0NuZcYf3VQaW67W3kQnWQE4NJc71QF8jABb
pOHoOQKEVmKoXSFL4juJZMVVbGGUWdEUf6uD0fJV1hSd4VCr7KseBVHqQBNX836JBUhF1Q0VPS/q
qEyi0Y7023UagWwy3iNFpLaThbuj5ua8EhE3InQPulYEymeGk0bKj7fjmz5fLaQxpDa7JII/INrY
cMsgv3n/XWRU2SUkvNfRvPWTS4J+5ekhschJFPGKFcZJ4NpNzeHZ2rNGvuCAZQqVM8GqetiYsz+b
pHzscuyn2jTKC4UaWsQUNqrx5rxeaYSIsI4Z898jMpzLKiGJcXE3j7USzi6JUoWqmdij6EJ5M/Kq
JFObYcDUHL0x54D8AMU6F8+CNbcKMMyYAtcjsvfaPV9qcBe2+qfwUWcpQ+3QIzEGNLrnDg+EIEec
o+GvfSbK02WkYw3amOSjyloUjNRe+wVHj03LbwlYuvJpVnz4kvoM/7l/1o6rxhhtyR2bbpyO5sQe
HiJIP2GrCIs092g4iDX/BWpcUt7pAKGu/MJyjfFE7SaGN6Z0EF2+LBFBdRXuRGg7vld1t+5Q
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
xI5rRsZ8D/mWscsXgMgqvONi1IR+WUmvlhOeHpoqbkmGbmmCKddy2Qan/TbchxUow2f4O04cfAEu
JYQ5L/DafoWEAHShGyHztGxj4EyJX7x8yqtcAWwgcJlMfy/2Z+sYHVx4ASnUNZeQ8HXpWibYIZuP
FjkTNuAr1SrdQnqwhH5cviaA/5OheQSigRQCP8RRQlRyBxc+biSsCZMpGISZFX2CZjSyU+7V2yWW
ay7r6zDWmMmDZjudTCI4MmCNXIWpp/bhBBuYrBSF+L/5EsYX/jb3bbE7tKSBxKDVS/NsrCqqNgPq
LE6lSb2eW+8BDcfgsBxnkhOXEUv0U/y1UADlGQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
kt+7rNkOSYrcXqbgq36Tjy1mVNbqyEaJJcQomY0hj5jTsV2loT+ykCqTokaSF04RFimKeTBrbOMs
fGmY0J0Y3FLdb9mRm02LfOxlSlD1IAUzPqmK1XSR8d/4MtempkKY0sPLjad2NV3YwFQOuIgbOEwQ
WJexgoWi794m/yDoUFziRVt8L8gAHObe8TsXdCCkIFw1w5BV4qiVphOfsBcAFfGjk1h0eqKL4hHd
+knMywKT44w7gE4DaneMKpcCfQ4X0hNR6jP67PdO/EqqXFjgnAn0wypmmiFT+lBYDb/eP0n/hSzE
W8aox1YjaQtyA9zwXG2XZMpfhHFKcSJlD/u2/Q==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=149328)
`pragma protect data_block
RvX6YNnGq/QfZrX3+SpkwDzMRMPNyB83XtyOs+h+gSiynn1XhUeSuYChhjzO2tVQ1rH3F/vCPrla
hD6VUALEq148nibJmMdYwv3hTk+sBmRcjCK49iKFYZ/tdhMSsIm1BIZrY8EQWICi7teBeErv3NJb
dWXAjbrToZfLhLs8dbOHQ5IeERmI2jxMHlIDLlxjLEHqV9ybINIEoYCUNFIKX8yrNAOSiB62AVk9
F65vgb+GThPHJp1sNpOWimfOv+/6Oo/W6BOOxzOHMKJY1us6t162gsKUU0fWBNrCj+vssOQq7SrB
crH9zn+iMCxEK0YZzuJkmCMWqZ7AZwtfRM+qEZNUA00xy4hADuAOa/xj7enRywhQzcafss6zoYIt
1lhyGaSALH9yhQlAkHYu1D0CdjsF2iZjIP5bXsPkxW9PLppuaiXqPlKiBsWHlmqTgUB8FnhBe7mM
kFq1zezqUIAflT+m33WmUalXKUHOqtdd0635eqO5k5eHI0wiUneaFAdCPFejIHyNFPCTvUsYCHSX
283+wbe1rbMZ+2ed6HIEA+kaaIKAxO0MLoXJGZKiTILw/G39+wS8OT5Xp5tAk5o2LnWbCSE+bBS2
gJ+5EK2PMHiPWhrKT6aXZzTlM7gHQn2cd7Jclduq5q3iY0AL5/AuDwITwSYQH0twu9KT9ez8D6tY
OTgXHwVBQVIcjZSk0pDezZfH41cqEAfu46BpbIxWq3h56AqwZ8x3EgOHLpvpSxxklNmRWyP2EywL
hh6m5Sfl84TE2Tr/AszoeaNR7okijFln5rsOGxKv+24JvMmMM0FSuhl2aSQBSIJPANY92jF+/+8b
d9vF8of5V+KIeaU7PAGqfuxhBlqWBQ4zcc1OvV3kUs3LxT1uBKtT3swa3Xja3JwFUolzJE/zx8cR
z7XR5sT319n6K4xUvhD2naLGMsQ5G4hHNsfQp2+wcSNfTtMsTxqiFGOaH+BX37mM5gnvUr51P0yb
yc/SNgXBvuBEoSNyNyGjUIFjxoLXekSooos7+DdzGJ8n/4NBrK693UFRjkeGOx3JDi5QqThVH8Kh
mJ3tELLl6f3MBhJcaaBUo9AHuCJyTtyLiS+i591GJajt24K1tilzt1/1PoF81irDg54UhB+6aJCG
fO4wGlJXfPVoFFbzGTjI4OU4gKQs0iLD7wQZ3GztTYB+E5MqY/ghXYQ3+u1AOPqv8e6cuGJI7m22
Qc+heGoOMGV1AIgCZFnNAOdnEXSoeS/QxnKGDaA8btg9SltrG/kVfInMjJkd3UvFpybzM8j9zs4i
gLSkVtdoByly+OKTzHRRPrDSoMtAVJ0JmXVgqkVqJjfy6DfDj5HrwLQQx9h5Kdfam4Va8FNYeMij
spsIKGWJ6RcKHZ40nDA+EXXhyD11fTbRhtOc0ui4+7EjzPQhuU/cMKeMSm7e+OFJ8LImQw+/Ufq8
qJL2dqTLUpgM7/BGpPcVIzj75dPF+fA9CELZ8hPE5l8i1ODEWil+6/rgkf7qIzUVCHt43ftXHjD1
F3Yns4n7pkm+hJ5xnBas7RRxixizD9P3kSWO5gTMuvlm4M/VjAtKqiQZQYjkFkTg+FG7I5rlSaIV
4Vj8GyaMp5l9TFTY1Bhl+pyN5PVzhqPDCh3Wd+SGQdgoGy9UKVGKnpGpt5978QaO6osIJpaAZ1Y9
h1qeOJ0WdB0RRjEEzTGaG1Wt1r9Rbzq3v9hMR4ILVkNqw4q+6krIiwTFgZvzRGjDf38b20MTirr3
R+dmuIMn9lgkadbWSBfV4mgsAUTCdbENmy1X1EMJLx9EqhCQkuCmCvZ89lAwfaDTIDmIc6oX/4Nl
UMAntgNyIF0s0IbrVO8xTbl4fSUohEGvrjpiUwcjgj1089urUr7Y0sCmZslzqBHwnKj8UQHp1PvQ
0D4AeMvJuSPOLCcI9r3UnwChSJ+JiiwfHwZLrlH1/hWe83+elsvPMuQp6Usw4HuRkAgKV+X2Peo/
p0N3EQaYbeTKu6usXYwNjwYFVExOeEFEglkhmFT39ArB4zweh3IhzbVfH5hVG57JUv1IlVHgqJ1i
GILU6iNao8AJRzB3Rdjh0MzFVsRaIPGwZ/P+pJMAaLFnxYVthpP9RgEl3/zIdDsyl5v1iWta6brM
sciKYIDuLPBH/hEI3RFwjFSZBV+5vW3PgPDY9DBZjH/FkWm0FDxWfsgUiaUdEMB/mk5113EjRgua
dD+8erOdgkK5E0zKrSO3c2qW9THrbhqL9LDQLLwzki8sWQY8IBvqvfU5ZK3VuJatFwFJamv50lEg
A/5tOM4vLCVq7Uioy1VjGNVG74uyMDU6vplCtNvj6r/9tLliEoD03dpoyeGp4URJoP+D38c/k3Lf
TgquqC/Vv4+3uugECDUb2oqUN3WoG8YEFq2q8xRIpXaSnzFapG8ygKqK/Lzdq16GOi8aJ+AXxlZ0
yHtHBBVt0t26tfGB3tz81kFRL5r1lpIEDsa37FHzOU0x+TMoZE+9EfEaQ74IYmcB22cF/AxD2ACV
W5LqvppKhDWzBDfOAjIY9vi/p+3rNRdq8BnfuP+33O2bQ1ZOa9FMmfoV95DmsnzjNyXrAvmdLBMe
DjZTBuW+ZWPZdqbug7zqveCmyamASgjP/uEiPmiUjHvyU+JYh5rXqwHDYglUNfalNetTq7uIIDF9
dTMW31JA/nwGhRKIUlyObCSkZA5Hbtt6JxHnWzlMicupJgDjhJcYkGrXBzp/q9UuUtipD0ip7c6W
iu7I9KTfY4qmsvTzu9CZ8PcP1SAPCtSoRxi182oEOrg2E+4TZDQEZV5qSAqqCawTzH+zXCqteVi2
YdjewlgPczPm80u2AIPdcillyGhcUtg69ZU/9/wYpH+EhTGnk5+GPBak2mcQz3F/PYzGAULOzSRW
1/3jJ/24NYrLrmA+gq0gycarfjWhV7Sh1WlY8mdzhfobuTSXuiQqHZT+AJ309ux34qnfzQBpFos2
pKa0BlyAZkYoa1VAHSsqm7szVIzoxAfxJ5T32rRcceXfUF1wWS0MUx7Gr2kPkKZ2lcjw9b3J6Km8
l/hk6itp5RQV0H2ssf11TT9T27iK5s99bgIjwME15pn+CIhLhBWdAWzGdbkwrgkHzisK24PdcjAj
4aMui8ysmcTvy/eAeukI6QfxX66tfzeXymoyvrzrJ5F3h9U/IY+GhZSiTot1AFKWbV5vFRAN1YKB
8EfKAJkgD2SFoTYY66I/GpT4QKXQocVu74Ju95lN7U3ffrnqwykp8I1q2WrB3D16vrm8ublCOtmf
j6G1/RpR0UfRT+g8DqADNdpKbCokIDfi/I8GbQr0wh7zpnfexrzYGsq+haweGyrQuLNjH1+BOMyZ
YBPH4RPJAXUial8A5lDCtd3HuVrenZoOBFxA50RRSHIJK5ESag+iUgsBxqhgcLtYsXF1W+8lxKsX
1EPGK6JOl65DVS0/bj4MDOVxC8cNgB6xovJgN/+Zx2qJMu7inw7hXSmck/b2y4HGiX27CJXFZtN/
xMF3qUw7y+Mk+w8Lr26zk8BJ35YJBArrzxT+cB4mGlH+5eRp/AMVN3GoUd+22t2WvMYZFqk2bo+R
dIIbYmtDc+xVCstgDmtIQxkI8YtqWby2NveT5CQbi5hpSaT/vAfdsJeyPh9jZ74ZI47cRL1YVLyK
4i3uxjzoqNcu80wzn5+NBlbHAdd5HTQVAc4NFkeqWwUcYXSeC6hSfUmBqdol02EcK9vemvZ3wbs8
Et2F3WGfPCKCJaT1bmt/9AApIYZjWMu7JGoSZP83u8Y6fTNOPOvHSZMT5SjrmLPkOq9AGzZhkIM/
wTpGgCQLIw8wIi3P3aEi+PZ6NZa6R9MvBWqoDxkC7JAZ2nrJpcBSv9F0OGjPpjDB9OE1L9c+vHWD
AvufAyXIF8MA1pME6NB2VLxhm2xAfGP6qsNDbvpjyOF+SKS8yDnePIsAepgAUScpYUKsqll4Tjl1
3GiTI/3qh48vNaUJDaKwBRnejdsG2MecuX40eem0cTFMJ1Aoqpqas2Ypk1+U3jBYsyKNiTbInfDV
tOoehBOApZWK26ZaIuxIfFCsO2lLukUqM36XCfaMvK0r1uk0tP2gfpDT/9lf2bK4xCVjYs27/V47
sOTaiRGprjfwjFCG463XdK2fsZTXvvN2mmTWCqRUQTejn+2Khhq1k5CE2kBlDI4u/ACfDDb2NW8G
TVA9yj+EbjhJ3GDS+Jx9PEI9z7ANQf68g9euFVBUjJUBKYtOOsCa0FR/j6ax2psjS49DxZiQD4Gi
Wie/HeOfC50J/HviJTkzEdwobpI8BS9jiiONu05qZKMi78NjomdzG0+FViurKtgnJLTk6Ei3Izah
2VCNbgUsQEg1ZUL20uIs9ZQDO3ZAtWVGgQxou1umq9i2iL+6VzXsJCXalKjaYtrdjMgylQ60DeKY
FVQGRcAZTIYmAeWDPbQSkwfCoS0hFE6mEecuR6rrJs8pR4g4Kv9GSTldwZMzyd20IqCZb8rCCPwJ
nJI3IBzQtqgcbJSCBliC9tnQK2ZvJLrj3ydVVbEnxOBDxPi0JV3zzZ0EEEDdnzz9sie4m3bINQnS
x1jSELpKfKt72XM47ZoBcrHga6y8PsVRoDYlYaZbBEw/K5E7aFzklQGYCrfDkwdk1NDd6dYxzSXg
5v7MugZv8tYFhr+IlhoKX/MikL8146TrjAKk4ZD2u9sbay9mVO+T46sAHEaqy7ZSV6WtsczMAovN
rILMgccG00ssU4hTo5An/hJeE8yh8BrXTZ9R17DDqSOBAh22qkMtEyBeL0gAopF3vuRYceD6I64n
oxjk+N3zEJhHvpcXItO2tneAXoGe+QhbHkTdWsznTh18Mf1sVv17tXwZ2s1S3DvFjGDYLWfufdPt
nC4WF2oG+HoTpzSD4GV8w7DUL6o2yRIPDRITW6fvrsRr0R0rC9Bj7AW2lHkWgrydwKILe/7Yro8b
tJ318zUS3n6Glp8HOkhlPgU04UyYo8/FkS986X5JVNyld0OHSoFRyp/gfdsFLyNChhCfNBXqY+lM
eBS5Wv2bdsR31nBi8lIpcM+pVmvlKnIwqCf4pCKJy+vjuQ0nuL5fFCCd9n4l4MVoVdn6HB4vR7MI
3CP8KDpLQiND4QBU2/5DQA0+vJfKxj5wLkKXPdxvu62d+uddmk4iPKGY8fA2QYUp4ikPlQm8O8nG
hTN3PEdWcbSiZgVzOOzdW/nmTIhtn0908oCBQDF5iNydGrDtTD94OXw20ZScCha6D/YrcBVfWAgH
SjSoMHPzYXECVciVox22Tij51e+uhYSnZKqf8gYZkjJyWC6CHUvGr2Gt867lfDEB5Ebjn3aTWU4l
1NwbZHj5vzSEqDOwxJHMgeTCfnVYaPgwcGs3/q6BQx1sgRSQPuBMP3sk3wisoQGUyoTyOlpWsOi6
faTVHqoQN76liBw9u+Kk3WveqqI8A0pRalWEJqseTiI8BlNJRWQE0+tOJCHKEHwFf+1flHvTp5by
rS8Y47ONFDd92byszKG6TB4hANWUhsYiph8Jqo5Kz/bf4/gl8m6Ujr9bx1RfDpPRfX3HgRSgAh1W
zdEe/+BjKV7r4xHXdaYrIfgpWFLW6LuZ807bXnskAbhXP0LjkubtaByv/5Ms7qssEYuXp50p72UY
xqMBIVk7l3tDl9V4Xk/OdUzXXevPKJdOK+xcuzydozjZ5S5o7Yy3A0kDkb6soZPTpHYjXLoBbF/m
di1SL6cEZZETNwikd5p6GbtcVvHGqxSZQ+SPmX/gzshmYp2n+r7qpEv2OCUAb4x+8miJsBIKk5Vm
VSLL4HibR2mDWf4g12A5Ay5FxpsDxvY94i75QB6VoS2wKyU55xI6v7f8+j0vGTcSqPwqjNMFoa5g
Mp6ydu+3TanL+TrCSGl7QuaWY1sZgCFWVBkV+Y4qgFD3439Bha5facmnFZsjxANZMabRMDfKGGMJ
D8E9VZsJXPw3bqsBwAeqxKtuZ7aTdk+YOizU/lel2TmXAeNem3GAmNBOWkcoirZ6IeKV8O5u104H
sb+wbnc/VlTnsPo6tVRcNW6I7ltY6OrF5kJEiMs1lXmoGv2gjuhmUDUhnrOsQfGexdNINBRDsh5n
P6f6PWUqS2Dto8FHZkgSCa89m4zggBGFDuhphYhvS8wUZact7ieBhnylHiw1SUp614GEtEh5DOTl
fzvSQRkiHZKaI1vV5gy8B7/0AkJk3mrNN9SDQsAyw5eaH7fWM/4Ix+QRCQjP8tg7HIDywvUEYpq5
pTfS1jjWG0XmuFkDzQ7kcLHfMlHDXN00xYwkfNvEKFYG8d8K9q1Zy1RDvZV2RxYGqN5wTVfy8nRc
fy0+pEFc5RQsaxRoOkgNOGMuM59JpV2aY4w4BWUUk5qmM4RRz6jMxxP6DZAWkWkU2hyNy6mDocyQ
g3mKp+f6PC73xnNrGuOXy0ci4Yf2UP9zHd2cFOf+Cw96aWm1ZlwJs2zS6Hms1fW5mRBsZcaCFsH/
FYjGf/XrRJKkLO58Muv9NUvjMbZhQcIvanNLIu1J4FXMFNcySnxTv7t9fjFG+x7iBftkuLiAdW1V
qFksZqgA1bVceEGRUDqZEP0ajqQIcHRwmvMG1gtSskrOS6pRAMKzIf43NPM1A8+R3LzDdO3+CX1s
Qz7CjxPg5kC0MRdlnc43HSuwzrySeye8QP0hy5TMB25DE3hgMNGXPvd+8c0K51AlS5B9xEwAgY91
xAgerElOaOWISGU7kA8pUyVZDAxJ+vlu7ccfLoEyDcPhLG/Ad+BwhJy+rmIuNzxhHKx3VTCtCp+b
d+whutMCcYyS8uPfuRpqxoEWOLEaHn8amg++R3sgvWOugNH+9Dyd5QElZScP+B2W9G4EBooCOtKp
1vQLPqMP5yLWOn9TvMW4zAobcrW7LwrlOrICpua9LEeyX9EqCGbcvw5Hvay2LltcAhRe95Q3hVzG
9jhOCRETOpxOix7KCOUSSxKpI6HXggSrcMcbU4RvpGWDMOGbwtC/UdwcGXuX50oTSGCqs+eEZ5oe
t49WtvE1JJyYxZ5qItj/kTvyLeysE5WcbY0rJh4zCMk1TKRsLGajspvOtYBLlsM+Hrqb41dDsfXs
9JvAxKbX696HibiA7f0t/SP/S8Et16LPs2ZQtMR4Yf5L5VsmavO/q4vj8fQc8XZzzDrevKrdbdEg
MMgiHrzI+IkaJXPj9N96M4nCkj2WFeP3oaXlUpjMXmDchvAgiz34zzByYTuwjslRQGPdo+1R7x5+
X64Vp2eZnAc8WN1A/iqGqDtKnWS4qeHgYrQ8TAdjOIb8FYJZaFH1HBrPwTT3Ea/AEIoBGWi4ieTv
B2rI6l8eQi8NoY8QJ4g66iyfP2HqLreCwZrCBztXZCPFKVbV0FTadeK8qWNfNpp5o1NgV77GU+Ii
LMldJ9Hg0Ui+3/qXj3ScaYVBG0Qt+XJHKGO8Va26W4ZH0zNm1KyAgLHREnT70/FEi3IayltYbBFd
0Uw9xuQMbeBdGOFgcnQbHp0h3hyDvS74uDm3bCutCiI3TBKoht5YxFYSlubQzh+U5Mle7MVpDTM9
tzGcz0UrduTKIUWpFBtdy5+Zb5qGvyA59akVbqDcCasm68pC1YUycpzVwGugDwXyu4mHknwoLvXA
7eyL6qAI/ZQdIfXLan9vR0wDwwJuwEinQSOWgC+qx1NTqrudYIauAFAntINTam2XaY0oO54LGIJF
sf2jmBMFvCAO5JI/S1oW2mlFhsvLkd/KqTDyPGHt49rWXRNFChIrjHhu6YhJbPPj7HQ7FUcJayq6
zJS2h87FTtSPxEUbd0a67dvuUrZMjT3/JIn0bAChWcPsYCRILz8Mjl2EKRHMvj/327FBGGdy54xj
xJEvKgbkToV2NdMj7gLFXbcTEkBvfcOVEdOVPyy3rx6zI1lx+HVetR4SfxLVKFrPg3mQ1fnsvbTU
QqtFoMC/2DPSxasfaH/UHwgwBDlLIS4DAmLwwnmQDWiZXLpNxlwNXo9AjqLCUK+0r7w9BaWF6fWq
tSaJ2BkWvVTXZM9AUBGU9540kRvaM9lv8Vn2W3hs828Gxvvv6DyVlTgoPQqftEGCW1EI3AjNlz4M
8QQZcf7V1RRYVILVQCccFQ6ZezozgII9SSpNj+CCQLPsREZpCV0lRCwNWMi2Kk955vy9EOqd8Zdw
yBfzUowzTJk0yTurKO3Kl22Bwya7GtlOnfD2aUJ7/gZIBexhsCGccg2n03WI/vCPopHkIXZ3sITB
THyJsxiFmIuNADMEgN9PeTFlJq8R0aOwEKKvvf1xWK4hc8YTbMBFTMrHSCLK4+zZdu1aYROqiffG
C9ieyrsjq5ZRcEmvDy5m/63BDdYvGant8yZn95qXxxuvuizzAYEKl3MsdSKp9mlvMYCxedocmBni
5tl6d7W1LUJ9L7Ofd/5EsirdAk+mwyVVIKwkS4rOPjfna74qwGTK98DTciXPtnO+QYz1uqkREvgp
p1sI6I86UdKEAKYH+QWMRA6OIZVpK6fr/Gl2VO4PC6q0j/nm2Ph3mwdF9qrJgzf+E4jrJv0978fD
LHQKPsf1G/q62vsBbZX8u6rOp0cz4bzLbeCaCvWmxTnUfbvbc37Z5vVC9DO6CcHjDSjtKWTpPAad
CIE/KNAkgv+DQfkBFNh9t6IUlEvtrCKutojZIbrXZmnIyZ4BTVDZhT8/SqybFz/qUojvbJulow81
CBtjHCTfZcWjon81HbK7r6NYbWnorOd3QE2NM44ett6oEauvywE2UmnsBrwHugYm5jd5m63BsfMo
uK4mMuUaL5WfEEwYsa2DNebvwPzHTt5uBFayL4ALreMTXhqSaVKn9LRvDtOmYcQ4ISaXHY42gzyX
kCDKTqClzreJldJW7Qn4ybKHVBtNTiH3pmmysrCf+fDr+OzwmqYzz2htVYBaIQ9/0kAWF9HN6asf
0HClI/YKgh8LPyJ2djDZlwwwp2JKC2EihEKIBbxJCmFOgemzkdTa0GJTSZVl70JWRNJCuqs9Xxji
Ptam1+Cd4oaQgu/5MrRfEgNtwGG5f8S63P5v6Iybcpog3S0Pafpd1VpKwANxy07hCdK9hB6/BGqZ
KpRCnQ8w2aoxm+KvSFhSBaFSP1p7dE1Yfm1THtZwykPGGZHSd16y8AUKJA0j1ra+yCmSHxM1VXcI
D+CcTfe50ThUI6NurxYk0GC2+0oqhHD3l1IQolbmH3kSnZIV7UrPlHK6SMtfomP9K3fXMRQx74Gd
RWrV2Sc6HKdAAvqHSYCu2DoWFptAgo+WNa+jZBNOqJwLc2Fzf0OaqzncsxgosIUKBxLeastxXSac
28mw1ovWE/N+oWxbrqXBh6YjlDOuMUspGxEqur8/W7aNbGGEHsfsV3k503wE3LaioiJp/H9bhkz5
iB3BUXJWK6HjVQ7GwCmYHCHKmGR4ZxRrbHDpTi0h+pJLXdwUdYpxFaqJtc461kvOYmdMb7nuDd6c
WwCO19hgNGEb+JCvAbuBr1wNNU5u4TUGBtwHoUX64e2SoSUz+ZE9zJmTMvOVbIdKfLjilPLhsbC2
6vIGFVzkuFf38MU/hO58iiPSUhCwSG61OnGNX8SPjMoSNk6IK8SpXenDdD8DUnXj4edMgWpDMGnE
O9hG1UUY3MVXb11lX01iSkaECg0c7WdbM6fbc9WTuyQPPO8hyQLaw9GRA090ObJehFfPy+OAcMA6
d4VBnv7B54uF9mWDcv9AWauvnq32ZWvdqfmPE8JcgR0//QLXGYISqIAzXmhz2xrccvbglGUmJVbB
ix/ty+oUQ3CG+Aw38MgqUNkqgUTinFY5XrB542QsmuMMmmiEDO/bpHGznTLePczRdnw1Mf7ZBIvn
/lgwSlL0Y6VPnELHJzkQONuMMnur2fQEXOBFo1pPOYDfUMVAe2OGAE0efkJiw9w23Q7fM24pASQW
sWfh5jK1iC7M3oILl2eEeyOKV31/zBx9KuN0/Qmj6a9ojm7UGqmpXYaKRazi9tJG1+9ojb6ykvIy
zbvEVnr9KdiEMGcSQ9sWUTs+6oELBjWySushUCNNls/HYGHO26CHcAKf4CdgMgXYP0wi7/qzTFgl
sswIETTc4mW6hp9PA7fjmu0BVR8HGBKclanLW947LxJf0gLWdbn6qWLHR/PCZkahEYzizulDA6ne
R94bg9hX32X69NryKEbAwO1mf6RpdJrR+GfvjEsVGA93W6Sba5RelaLVYJJ0k0P1pc8e+o2TwKwV
/tG5fnFvGc9FNbGTmPQipUOreQ0aczuwNVqLziiHIMJGl6Fp1XPon8TG3MH532mRdClCqzYDvyDt
36/MW+X8U6I3z4z+s3QK3FolV96b+YWFZcnpkXqlx3ZIWe3+U4scD+Jf4jdDUSZuF+yvll37ANjQ
ol+HFOZ+KgzVxxUS2FTdxx3OeERAcWiuSSsSRGNcbrz88S9GJXWVbNnRuQ++zHkADLzoWoyF4yu1
Xt7qvKpT/QnFEhXm4MaYqubfpbkbSZYMi2L+Du93cfdFIDXmx0DyTAK3h8wNh+SeMtm+0mqMj5t4
4HNhsjUqs4E6nuuR5uheSXoOKSv2Uf9toc3O3BScrDU1s5+4xsoT8ESprE3EDEvHL9wNweyy9It6
K0IPCYifFRRC94eKZeF379/89uPX5nFxAbggPfHCpWyrn8I+B7RcigBmfghJRRvxFKdAwzPBwWv1
6/gsvRCgvXDm4PXhUcNjH2llqgM+Ux8ydGKkBli27pQkDqStezVKWhBgCVFovI/DbaMWtWpmqgNB
gtyAp4BwFRqtCBqHhSu+in78J4NH1XVJWNj6hx6bMI8R9yAAYhA5vE60+uxOAxJVqIfmDY3amvJs
fplqjNPXnBeW4rvNvkAJ0Dgq57yrXMbsKdR8lVxffAxnNsDN7fOEjfZM65lG+h2eJ9IB8RwTgTxQ
iWdlosvLSp7GQm/Wh2Y7CCp9zFNQARbgLC9BDjvS/koGdA1Ew0qZ8WBqF9ikn8eiHJtcxgQFmbDp
5h8LIdvmCAVhkYYinJ+wOeq1NpVZIx6BpAIVWYQe5wuU+5B2rAFhOLtxwhmxiIJ7aVO0glTWvOnm
yGeeAqgbEyKXnC01iFg+Y+Er8LYZVKygOoUWc8jHRCD/dHB2tFKZk5ZnhG4foNVq7feyz2zqxPTR
UcoOiFii5FRojKnanK/4/NI2Lux+ECOh+ZVH3JWFYZjRZ5A5WIbktWzeQXLn5CvALKjDAXmMXRCM
7wd4kdRRJzuhdD3lY6HdRPhFRlr60ZjZ9M3smdbNEh+2mhIXJVEkYWGAE8JnCnr+TXQ4Dw/wjCtv
NEYCne/ub5gK29NLCZP8f8pP5uTH3qAGi1YItMXPwTFarfmrzdvNLPAmhwNXerjilH9ljXlw8Ltw
LB/2Z1X5CeK1O1v2UKU+YTuNboir5ZC1a1FIhpVk42rFqNUMovUkhv5H0+TWWsQOs/ewvXjw3yPn
R5Wm631SnUXaaImybC13GRs73JACoLRyoxCoc5v8MDMNOXIc608v48pS0aYfub1dxtkRFIily6jQ
3/LQkyo7xPg+2E777MKf++RYTiUNuGQRGK2TV88WUdN18SAK/uiS4Ya1xszFg1KL+AU9zb+tBhd+
hwnuxAuUoIjwEyZdk1RlX44nbCOySEEUHZvFVmGDowctDp7eAxvD5WRxDPliTZMIKGm0I0W0+pAz
hxUHR6GA5G7XitrDgjoxEe7BKhjZ/vAI2V6/C9nqJSN/CMs57kdV9cLR6G3+XANZMH5Wx3DdCBRJ
LzC6ZhL9PMiWy0hL7UY5Y1DB+zHqvpJfDkUbR5yFhDHO6kh1h0zGZ7tmiCFzc8LUFp4FdbrOlbIA
3rqBjoX9u+frq66Tf7dQR7gC99CZzxfVRkDijh4CBAWzFBGeqhetuzLqWICVGMTlb/ukO66LA03f
qiho2ow/d9Y11wh+gLdiWkov/anuenJ69rClpwq/BRDhDkbykavgzjPmSpjRWYLxR5doeH/HXDTt
Nf1fihQrOZfNJljdf505X7bVaaRpnTtlJ+6sgtje4LN2HfE2ixCt3fHE9N0KI5d+iwqbARUanF5I
1pWfnx7oS2rWClvcb6laJchV0P2YOuNm3PzITJqQZZSDqKhrgN5lj5s2acZp8WkyJYIDVGRP8Zle
nePDoNUbnocKpprJG54oJxc3Ku40PMlpieE/pdnBoHmu2Inn0KPhnyp4JyCO++JgpNBFIa2gWXkL
3dNo2g/BA4wItQf3AEx+FBLE7s0pIYo6IHy5B2+GzdiERmdtVTrT+QQIwXWpiCU9jROL/ijb2bbA
TvfwvGoaldBWyBefmcoO14HGV4rnq5bPOqeGU1nS63pbn4kezykOkywWFvkYgpW7Lv7LwetXIMnC
arfN4rwX0iucCWwCY1YxQvcYL/Q8cujrBy4s2d58iy4Jr+63eCzf3dvovVnVnrc7vkGzn54f/lYu
CBocUNHXgKpdEL0+yBqKBk6Yf7BP/GyDuW20lsjibEoYMyfgQ1bckqf2LJNcv+UYcxSEgZtblEKz
+VBT+T1mt+/O1F3vP0wLGX6zb/fCh+45ZMXZZNghvK04VgaMh8KkIng7ynX5M3q1wmzlBXV/vrmG
x0nXiMZobxOfaMjLzcPgmoDmTpQvIGIB4XEJx9DdHUZ6t8V69qHatqxja4GhS5kmlBH4uUbzV0BB
mATR7z3hU2Wqr54okGqyd6hsdiEPCJ1QV5sXR/Htz+JIp4opcQUjM82ak2GWU9cBuq9TwQ7eIK3Q
+KoLmZYKprD+UAD3ktzOy4QbhwAwxJ3ODZGJ9FZY+sQN7xfMMWH/C6IAz62ESS1JJvuoxFnhNzW0
sWPHiurV1uM38nXQJCOyPAm6QuU5v+7htmEMFCA24ZtUqcAil8kdEyDei51P7ZVG7ahPEsznbBlj
XiMVBrlqjBACUHWDGHgIRI/vBqDQWbiifhkGSTllOuldtmOex+4hZPJfhtekn7MAeX9lBGILW5PO
X/waBq8VCmDhen3KmIsYzvcuO2A9k2Vm1qWg3ZX1GLOJkFqwNBlBvf3QIi3dYwcRz48W/qLn+zQN
db8/72FED7BxeWziPUo9eobNO5Yc/MJym6pADGYNgZuAyGbs/2nwIvJO59qNGlM/VKUplLn6plqQ
Wt25o7ZEKjtyl2mM9CPS2gT180pyc17IW8iz25BAbJEzdVvXjGvq4m29eCKdqObN/+xEqiSWkNSe
x9cn3SEZgf6ZyVWXJjKSf73KAvjdH+L09hBEyN+zaNQmdqD8+ecaDwDV3vne9OOqlPah+nnU7YwC
2ANvcU3n03E1EJhnO3pkAYyJ1/H9wdgPHlvY4T/Ff8NdDccLLtmSHlPRVoHA+2rRijyhghHi3sEV
CbZQhtUdHyFCPfpZKmc84l8aYJOgXir/cNZYSiZmz/h6Asm9YvY28saMBZbI24zWc+hj3trBgnBB
MlolALzH5BMFEQQpQCppU5N/ec8V5YzVfmVhcKxlPZRlA23irFv+6eq9mF+cNEgfw6SyBJM5O6zr
3WjRfEhd6MXwIFFaFGUnT6IQTnI4g2IE86VEiFQ1otH+RqJtu+EwUzuo4t6nyea9bm0f19RvCo99
bXwXezLF2N+L1UM76g5Vc4evFKn1/gv/vI0g+y0b1qjLKsULuK/a/cKsUKgcaqL9NRxcoX+IOfpW
pag1VmoIJkHMgBjKBFJeVBg72SEmwvKDRZyG+nYE6Vkz2VdebTBHjPkTHr51Fy7k+H23RJh8ei5E
rHeKmY881ZedkykidsBC7Ywd7Mnf2tt4EuU/cVCqTocinin7J2XOAXCLiSU1zdBFFLMIgR1N/GQ5
PphpV5MJ0KmO1F+qHuO1QKWjqFnxude6N2+UklPcTDq8co/RlYD13pmTRgOQOotFQvJ1SmIfYd4g
E/IjukS/c97gFuxwh8ATJwZ32ZeL3vrGNU+uUGsCcv1TBovAHFr4rFvAUBNaTHojIxmn7+1S0Bzv
CVLqZ1bb+AZ6smzJmgKM9XgBdvXiakkFym0PEDY9L4Xf3YDKrUMiihejtcIBXuwX0M4Xt7W3tgqQ
cwWOcFIC7C+CHqs+QT7Z/zpW/rYa1wxCt6r6zs+WM+YpXB8fRuRJHDmreMFV9h4OxL5M3nplYmcV
jAIzbTfkYA420oygS3x6eD+/xdDZ9x/faN2AH/ayvy+ds7essNHnyVQyx/6ED0cTopHLH5HV/fBt
cdhtCcsafnLbcmdzXvbn15g9dn1gjP1JMAj7NtafenwUt/HIljOJVhCN3YeLjn6YvWxDadAQhQyH
uvjEgWERBPmwH3OuTPzq9svI5ZkppfdOfHyYJaPLWQoq3eL2BpAxgMHf4V+mN+WjHw6Fq58eBLDa
qEpDLN5ks4Jug2zhGEtP7WhWjHKw030782PEH8oEaaMIrcyTRC8f/G9O8TbZDCYWdTE+wKtNCHPT
K/eEYbG8u/deBSHNUzilbid1JP2WR+rclX8TpmwEIbujp32TBnqt0fEovxJPr+lyA+MijWtPf9h8
YBEFXXWUno26HvZ07g9Xu5rURbleqbyltHL4ij9ER8TjFOtEp7mBt9XU7dcZ1bUjYCJxwX9sa80B
18aCRfttHY7dHL+8S8w8LQqlZkbqhwG9CzIxGF8Jmf8AmovRUNz3pI3VNBk/IaKS8nFjxQj2yDJ5
ThPP7ydgnrpBGaBYbGSVjQmxEyzlp7qTG00LqTdTuo0SsrQJ4lxyK/6g4dUhwspcgD8tEA8STtQB
p78o6YYvpH8ARFt+y6kCNdWqFyZoYpVDSQOLDTtwvNxAXQhNGEoAHosDwv41a8xj8nFTNiECv1am
3OGI3L/qfQYormn5tlfL+04unSiCbEIFwyj3oj1jSeyDCiWtn8iA2lVdDFiH505P97h7QY2rhvAi
Vp6kleuRST7Dz9xUoHWItyMZBr61rC/qhFh4cOh6QemzS0DouT2/15ZGjrv9WAllW6tK438VXzoU
2aVGTUxvBEKwuazPI99zmY0Gd7NSBEigKmkvadZHQn3c0A3clBemEu8Z2hwYksm6uSqga/xjd5ii
BKlggcsjOWrIAw/5mxK4vKfrYCUb2oYsOor0HIoGXIBT45KqMRdEIN27Vk7iOmYUoZHfQcZ3SYiU
5hUiBl8DpCp6VAeZqB5CvmztCMl/EWYuMqy1iIbEVcyKoKXfm2gKh/vaFpkdUXUoy9hfNp86XgFK
z2JRFUVKe0na3rPuee2Qyxd1BN/0vToMqLBppDBXithx27HeNsYnRhSFnSTu9pyGZAgaTeiZ/OAv
FjYFITwXbS6FioRPavkrOxXymQvT2noiRwK2Po/LLL2/8aypC0ZT2J5fGsgpnVuEPTQeO8uns8po
C7eJFvVYqSwBXXhEuBPSU/8SMFU7d+sGXHGJ34TDd+cmrDVNkfQl027bQX9PLRAQ1WUySyYlIKJv
M7z5X7fme+IJWtm8kgCtH4mkwSsjGF+BylPjFsB7GDP2h3rl6pWCRfHP2vfENkTEOWDj6A3yXmF2
Y4HCXq9LQdFGNLRbsgw+SH0Nac/N/W7BN1LTDCLn2MCTKuOUAM8IC1iwSsB2D4/YpEUZaZemLf5h
CWeKVqW0M+GZUChhUIr8lWCkFxCDy9TtsIN7+Tkoq42P/1DsnN+IS4ahcmFfrEnN1I8oYDVBjg7h
AtmaAbdqzvmsQeTO2vhw0STCUIOEVWpopJqEZkc3pHbRf7nmoHfEE1hQ58WEHSCnIF/9WMH9XhPO
0O8s7F0tEKAm67pwgKXlSyhwJRkzUZUHUu3n0JXfeUdEP0VnqO1+KN7u1iPEHP07/0ZYzCl+VSWM
Vlk1M9RuknvyvCAWlt+pwOC0ggodtZhUuchUI1WojFVY6XxNQ1kce0yjIxbowI5sGCxzS/UH6UII
hHAnCRLE3F0oEnnu0rq+xLVdwnqsG32T1qpOcFwHi/K/6bTm9UrSdhFdt7WhdWr8jA7Vd4ETtK4a
VQDW0lRQ6RBhn9yl360zwPsPaKH0gle0TgKr1/fhZ6aaQNZf1Kj5nd1kujbfWeVmbqxSnHZu95Zx
dhve81M7Y0yrmKTcbpmUzqKiCCAdWjA8uEA+sJD/Wuq1rVuxexmHcKYUDmHm4b3mbxD3ODRRcLZ+
aPK9ipkEtZHjxyPmkwsbO1Lp8CcVka33KCAAHAT2RGznXSaVcYVDFpIw3tGrr6AIDQvkelJq8mxW
XTS0Y8CeaG7Idxq6kx4arJqPXnYxUc6u0K9yF0iC56BMTJxgoPaIM2PFTyEKSSiom6d9uQtSPyz5
2+i5lxFW1TkxpVOrtO+NAGF6s8VkU4riDvr585ZASSp1sK7a3aj6SFr3hTrDRglF3O4X62e2R4mC
Evsf4Us+kqou95tfN7cE/jLGUrHvaXGF1FsqCqJTY0gvqQgbfwdx2RN/BhdrUaFXAIsV7CSpyFuH
UX5anPr01h0M2rjG2eN/caV8od+1F9hcubI8ns1D9xVaPNkCXirKRsvQyFXq9g3OBQNWJnrcHKIN
NjE/qiLEX4egwTDjJN2mi0l+9OF5VgUemSKR36UKrBgK0QmU3fyRQhD53oKFuelmdOpUMrd8Vt1n
23bjuCIzN1r0aaUSP7HNKF+6agC/+SAWGdtIALthvk+PcxwNpfHYE0b9vbVJrzwAdLHGDoGe+k6q
ShzlM/2DIaUFD/lGervDeRVw+2Jdy3mFvg5GrCARe+mt8wN75UHpMTePYhXmqj4YURm90Trhjqru
fI4TwpFicbES1uUX0FkM+Clzv/2MmGVWH6x5hoaNA2Iie8NdHWjU1ZMQnwSf/W2PKhLUEpDhClmJ
kxq3cVRtexP8jWYTnMJiOG2Bl7/dK0Qa+3prU6AWWSuxcmLDn+tbFWe5IOlu9Q9eFoN1L1an7wPd
oMvs+mE41x1mclzpPVF2bSzAUzHLhdmIiCACuezOoi9++jw//RvPIFFpCv87x8LBzbOSyQwL8hSM
quW/v138O9cTFVrqB4oWJEAGkMZo3f52RRLKnTJvfb1F2cZnK/mmYXTXLMdIUjSODFFO+UCYhv/P
3twcp5m6wxCEg6hIuOhBK8EIaaZKtiM3TzJ8++olSwE0Hr7SUfze/7AOlsUBgMdw7lfUbCsxEH1e
ffSfskUbe0YfhPtA/xyqdL0cvEAeWl2xjdSCVwLPo9j7o64iVXryEFvu7DQkEyY2K2OG3ajFejsT
D+TOEyVFoW7vCdsceAYqTMiCncnB0s+hVkiLoNPVlGPshhhqbxvKMe8iS0m0WH3PIrn+1gnt4tlu
GFtUJ9KFi06usN9GAzbPkHjSZ+bvFCrtUYNYfkJGrc/5Ey0sKclor4/goAYrYxP7JGf96tyBhMOz
hKFqooy2DhepM66hs6Xw4hsO9gLDggqJ7bMPg/xZl0/hrKRTaYBjPyXnM47MMOejeSdz2h8BI0e/
HZysqt1VSL1qJqEqfoiStx7RHNRMImX6aRGiH9baqE7LLqfDbCXrwXmW2xHVj/R+lkI/RvsTeGZV
XpMCggZNwsRXSJmaVIs682sOVtjd+tol8ToNt/OURg0FehD3c009Xc1kDpNiS6Ag7MTChjX6MD+m
/hMlrqO3hHukRLhRN7/PmpG3yRDe6pO1xoiO9QniVUl4NyuO2WfuolI5aJp7alzM+fcMoPCi/TKu
wPqWBR4lZdU5ZE1lUJFSu7Zreywv+4Hn+ME9npR+SgT+xIGgdImjLMwhW6rXIhHlxBjfXyxenu+X
Z0jGS+6xKYjsoJBVbwmAXJzaN8zJ+U9Mhs1N31RTu6MwPtfFvX1Eebxue9/H2FZ1X4h3c+u2XxKP
3tkN4Ptexjyii19r7jF6E/rwNdqYP+UdekLK+nSIo231Ah6yQjPNTsOUjF3GM8U3jN8epQDOdJGV
T3qkTtDuHIfxms3Qhs5YuPcTLaZdZjixiyPb5DksHYcdopziaaqMll9c3qQzCo8DmwRaA0gFfxTT
hbFA/jjSSSSeGA6VRH3dFFNgrkuI3cv6wl0tvcTW0O/PkFBo4m/D+XarQ35xHzMmn/hqeBAXzm0g
bYOpVADvgzF5PKm4v7A7stPMgAGA0Z9LKmlCanbMPZU8JidCkLxElSuAvKGRbJhHuPULOBzLV0d6
E9vx0jd5CumcbEQ6z/4wSlpuAsSqhbPYjoTj4aH5I3Nnnx+wdL+8xtLwr/rkIvKZOqGllkC1+Olh
jIOiURmuaeFrECe3/KFu0anw3zg1icvfNQwf7SEPk4bIjTajWCaqjTKHolesW9aDJG3BpiiO9Lj1
KLD6KtHTATvXuITWTnoPrmcD6SzaGMO4q8qksgGZv5lliu5TDPLsQq+iRW1sr29ahAeThKqBQL0B
aPXjwMBqt2/oldHyIPASzlaox92/KUP10YH3qcTJkB9OeK2J9Wo7nTnuKpXx+FWSA7KIyWxKzc7P
Ywa0wc5ZMezHkUvmempOiMrhiXh684cDQvkAqB7++UC4d3qxruvkbVO8yBKWHFbjyB5TQUxZnU58
vRebaMMc1LZjh0m99n66u8QNmhTA+y7tWKMWL60xrMmR0lb4Kq7OPyRo9s0t0TGnb9NG0pIqzOxp
xGIqKVcRDqYZW4UPAPWTTXsmcY8SymkXB16zHoke8d6XBxlGhPk58rY7a9f80RkWg88eLHPZUF37
m0PmbZIrD5Emld0qYQaoncsPYX1OdknHx77jbpH6GCczA5ZxcDhKXVc2yX4TGNoHo6sM7mWBsFt0
hwjFibAs23yz8YLS3RRl+ehIZVwGYvIHHm59U6PUiBw0AHFh5VPGFaC2cEXPa5GVdj8gROAbEnMq
NcbsNDUEYaSg+1MBSplY5TV+rNJBFnqqRu61Br/X84W5xujgWYI/5rAaXF6RNblckoCnyhTPn335
y5+xgcAMLhgk4z8nNvkUOtbcIbtcYN0ub4X/63iBvAea8pOMT2G6D8KR+oe9Ai8urLTHhtCqUhVr
CCC6tSQleQKXuZq/G3TfQ58mHIpf+s1Q48g+evRayF7dWDjUrqEnxE0+xeUEKQeE6EmNcZez4NAJ
0N6AxM/2fBoCbK+RL9MgLp+IHKUUHkJ8Gr+AUn4Q1Bqs4L0g7qIV+xZJjZlFX3bCr8A3qBo+Vbaa
PR3L1Td6lyy2PF9oMHZU+tKsPTPa3eDgtXPAUTKhH2NZYWYvNi8uD7k36waWawBxaAKb9Q92Mn2m
Ck5UFTRw118EFv/xmrAE77kDPfHwnSMhmt5YR5J9hLB2xcS2Nm/IynWVcRX4MfOAeedeikya0quG
xJmSTY1gn9Q+E309mPmGjawAJXZMboDZoW/wpApbUbGkcyn2nQOwHPInPiJWm9kmeC8edVvKX1+4
JH1hGlJ91/xo8mwfjev0cZ5CsGSXTs/IuDKfBLYCfxNRMhSKoRiPgPbgUA/qA9PF3yXIpJ9kPN3L
U7TYtQCkTNSR3OojyrMxnDfQzqfNPqg5/iggjCcLO2WOQ6gW63iTKt+2eThtvG4UUavnwNhsgbZY
4vQFF+WtudJkCR/5ThnjO6vCgkrhwnjTJrJEA17B4iA9YYyVQR2Wsjng1dJY330B02hTkpib5IxG
C1exLpL2Tj61bRjaO9SF5ro3s32uCP7ftXMJQ/M9KqB5EmmvsYqVN+21vqeQXUIZ6eoNUtHNcucU
quxcH4fqfYhhSSn7vRG8jRORidGVX/dYOtgueowRo+ZSsMIqtGTHfYgNYplMzDxEEg6e0zFmbSlE
vKgA4/+y2PpsXl9nqV7WW1K4TYTiN+TY5uPq2PdIwt3pTZ/eSBzC0IwTtz64ZiXqCpFLhq6uKcI4
SDvH90ZSimSDEi/EaqmMzqFV5vYNJ6xZYABUvN0mdkWlU1mb3DvS1a2ZkCKaQRgDcwDB622/iFuP
w+TH2fD6/LCi2W8KFBgfcFXBdm+X/Xnq79cxjCS35Oz3bt3P2fpVxXy5Jefd7UZOAQYroLai/Rj/
8UpULd3A5ZNcf0jlrHnuB+jd1Mkz+ORufU06l+nBJQGS5GrIhLvAi8n7rTm38QXlJdv2M3iPQ2De
Q/CKWUkf148b9idMIZbiP7NYCpoa76G4jmzGTvJSU23Br9J+P4u+e6odDjcIpngrvZVhvjQXSF/G
lxFO90vIhfh+753TUmE5Dbb6wiopEzbR/yi/fws2/PRZzS7VwdY8ne+c7muvb5AV+W+pKxMYbJqp
Hw/0h/Pe2UgdoczQBRyEgURQEzcCJwStiiqf5FnRBH1eWPRGgoVoNSeVciPgspD+hU1jQ+r12bEx
9EnP0+WCVU+4Tck4bgt/GCTEYR4Ds3gcYZpCHnk9+PqxcrpThX2OVgmFxZtPvcK0cNVSo8ymKPgR
/ASC83eC+uBYNHx4CpxhYz5848fM0/EGaOHL0rdjN/ABYeQu87V9FCkvXPDkmrC0eqebFU1EkYsF
kSMCEaA0sWzlXwB2asIRhg4KJpKCc8WXIXl8vT6Ailnh9u2QJ60IXghPp6ylUo/AkSWmxOCu3aPU
29diDnZHGZ37k1B+ySnhpFoyeq1IRLNsqimGv3h+ejO0DyIixV3CjnPmmg3RGdwLs4/u2X++41oD
MjeaYEseQCiAQBulEf0qasWHE8P1X/5zcPYxJsA82/QjGTWdYnbD6PIbmLD1/v2EKfHWb+Ifa6d8
hMzTOTI/f8LjiT16byFrnRfPp5OzYFiYaoqoUeBGS3PA51Qd/M2CSoWxgrWn/ommK7LfwwFk1MZe
dFXRBwZILwX6/11Ho0u3NrcPVYVDWCZotD3iJXhr6Gu0/F/al8DF48fEDvGuQjeFyJHPNnWCS0jI
GagS3xnXCUUVxrNwKkHdJJvAIGnz4SPqYC0v2rnCclBQGopqvYuejhCWZ6IgjycASYs7Z3bLZu0b
xnr4NuZ416x/z+gQkMUKBfWzpaSojfTHSOMd9dG9qlk8NfWYOsJVBdlnVRjVi3//iTyrKl/3TsO6
4/atHu2p2cQVnFkgf2Xb4k7zRy2Yp6jJZ0Y0ZhK9Y09RCzSQKyzmGlqxf6YzZIKeV6xQCD3n3eR9
3qxCP7E/iNGaqkRgI/JhU3OEHM0yA2YPJcjiLTsw+G/KiTCn9CmcX64xIXPfGBl5rKMcrL4Glhl1
Gh53Ci2aHAT6h7B6iBuJNAF4gEd9bR7ZlsEFpD6c9ifGQ5QE4iQhsMNB47hT8J0MohPqaYCOtTYx
htCh8HpLfw/ikzPPIM8tG7tYsKErJFieZoxQBQ2TrTiCKfCpp4SsZkZcZ7oMmONMglpbhcv3d7WG
f2h9XUveu5jKnfo3jjUHOyWo8xKPYOGrjqUVbdNwGEQh4YH3+3VexmvdW8p7F8fUNCvV6hmbdiVc
GoxxFk24dGo1i1nCm0NKwg3AtIv8V+1cmMkHeNeZ2Ny4t3a0g1UYoq+0CYjwO7pYmMRo18gkurK0
W+UOI2rb8OpdhWzHW3/w/AaC6kDDzNEX0SylYJ/NBLp77Cmzl8TTN0KYJEmN8bxi74v2hpITYrwU
igOsZMRPxsblcNEWvHQjwfoEcCxCdvL/uIT6C8EJCxJOGYP+ndybRHAavcgIygNUCwa1Nk24iDIb
U8gZO5RrrylSEgNja8rcUsMcYWeC/XWYBPAAc4RZqMmlhL+pZ2RYBBAidfXsJSkGc/wvFAcB6ohM
u8mWL7Rgx0CmLw0E/IP6xG751HxsyLNNra6y2eSv2qycwiyyxvCwJG1jbV16oineI7i2qTPZy/u4
bCPxCyMcR/gv3qivj4TSEGnjrCjDJk2sV8TS5JLtDE7vmt/uNtp3rGQRAlm0R8y31up+lozYs07V
2LZbKT/qzWmEpcknf5qzLeNYaLHWL3wLiNP347udGJ10ynh++mRyFH0e0bs2bjtTkXPvweb4ij06
uo5mnjnN8xwAi+AmiiMQwSrqDZMaUpRlliMvFnA2rTLXD4KAYM969d7R5HFeoFkjgp5kl7zh4vqP
SMEb/85OH8qw6zZLnkr/3kOhAvLSJeMzln6oPfjEpFaM76Emk5wF08o5ebGhrrcZOC6CQDCggI0B
6K7c0lZ1d4PXDTfnBaNf/YOFzvlnvWEa5nQ98QlKPvrT/TaJPZSXfZ7eytfIIuZlZIKxcCWaAS1E
utuV3/GxjZPaLMqbfSTcOBpMHyIhJxOovolJ+NZhVwW57GVw4qBOW+GC+bTxpSYwLeNJMzvZWudR
g7P+GAAFm/JJ08awURla5nS57fQGcrAJ8qjyt2GmLMbKSIWQLg9k8L/6Ij/Nl8WRf8+AYVbZwRTr
uqSV40ZOH4Xw9OiiFlRyCTzAONXhewKP8PtjO/UFTVpBEwh7A3cj67tm0WO01VOxlseERNZIUoL1
T2NGI8jReMumPTQElikfDZu8rIeWALZcl6s5U3mGFZQgm66xiOAsDmG3bj2VaI2hx+u0MONk5Paz
N3Z8PDwSLay46I6YMjCtQRrNvm+BL3V5/thtZXuAy2BORPO6hOAjvMMOs76agcyXNgnEJppEbD3f
6X45DR5bGsv5ssx8mOLgvX4dghDYObFEpYvvJgAMJ7atSrLuCaXo+uhFSvQpoSUi+xZghy3I2U25
YWruiautYrH9IRl6VxQ9rP+T/zwtT/edLNkOWJMUj9wfMyX9iBY2+IfvzPVFE5XPvdok+w4J2R70
csDq4ENq0HXNvkfRD8Vt967mVeuTgGndrQEd2Bys3a/ie5IB39zG1Zrc/H+7HtR7gqu99w6neraS
gS6iLJ0NT3lufxw7o1j5Vw7sMCc1omMG1YKPvFsxOmtLvk61Dfzuox9PvN2ZTgrbWGp+HMSxG9OS
sLLVi5nI/OZ1gXrTV5Y2uMHMQ8gqGOy59vmkbfbGmqaNa7/4tn0lqdDwdJBJWIa2sTUcc67bYEOG
qIKrQZndJdLsyDzcXKBKuf86aI1B+64Pf3u8oYhUzrmzVH8h6lRaOLuT6QN3hcVhFKpq5si5cAG0
Rl1NWALYxIrFkbh1tOvHJiRlJC1b0kFVUrdiCfvAoYxeqpXo6WMAFJt8kDuu+WpnzEeU18MUn7We
oYxS5YxouZ3WxiQJVsoGFlH+SxOgumxxFludBW14niCJsn2R4Qp9ja0IH80G+kWv6xf88m/SERxe
nDZngZS3CnG9hb4hkfXC/kLeE9tIlo5nIpZR3BXdhv/xgqRps4l3qK1ihrMkG4rCdMdHjEQ9FWum
6eCRF8aFGC/1kQEhQxMwV/ZA8wV+zrjKwhP8FIz34A+JLrnAJ6Ch2URokJPpim5f0Sg2yyFDIpp2
8vD0G5Z02Gue2BoFScpEvK0sAK3s/WgGYEDv+75Lm9BSmkUk8o0fNxjc7lrYV6YzYVqZgkJCCs9I
BdJSy2LHOsOIrI4/yPcsROGyDJ/LsgkcwMfY+uH4ykTAu5T3t65RUt4uy7hWQuwA3yeKsShrb4nA
W46L/G0OUGPtHG5v34oWETSYnAZQT40gcbsily1kRUIyBx4nydjtstU0eASv6Q63adLXHmgpiUQO
JcAdLjzKuUJpoNePhM/mpFSJ3Oied4vhYcCY2NhI+8oEBLO6KofmhgKxOACE8xLpyhDVAHG6yA1y
7xYRCKOrWDAQUFORyePIcxSG+zzoD/9XBXVThfv781VoWLMSoj19b3VG1EVxrJpAJqjitz/YZ8FS
Q/thQ2jrxRNgUYb4mBSjP58bd6xXnQiJqFfgXx3Xbdt6JJBH6g9m5URipD/pPqiUMICYOWQgVaHn
XAiHWDO5IteN+GAtTM19b/Rqd2ZRN6b3u2/GvhldmwqFxCuFIRQs4oz83atsLccRSyzkgDTrlCca
kaetuFpMQzs7xwsN1saMdf0jCedkmMGvJQdf6vXtpX7g5fRE8rvFS7KYa8u3I8J4KRtDZd5FibzO
V+36wrUwEdKX7T612ft4V60WdJENkkNkbSCgS+O37rAgMYLdpEP06t3LFx9PYiKtBbUw30+gLIWn
aWJBqJMrdWimVAKcTb2hpxSwlwXR6IAYiYW5Vm5ygFR11jfIGycoZo0+nfL8G8N45g7zYQ9EnK9G
ZYE72OF9DxZ2eyQDWseqh3Aj4aQkAaTwyCxkEh5TlrkwizovaSGxA58aWEWt7O4RvOIQhNp0OLrl
udjsl5bY+Il4ipNRdhLXDZTbi5LaqWT6pKWvOY4uE++ZkQDvpmv+1eYsVDFd5edwNovyoqTK8aS9
eJl0WfIetm9UFlXl7nOed6qOPnEf8vE/HfzZrKZlfreOnUZrkokYczfFkAOyv+uhau5tFSkusQtw
AIYWLhw+V4qYy/ZaIBxUpfxGxgEMkdFHeIinqgLkWsdA4E6eO9UopxQb/YI/BkwjoXuWzTDnes+a
haOBxDjbQ9ckZ9irjEs+NlFMfPWZ5798MLvzhn2sVUOrckXWwD7zCMOeT7jjNeTnDMtktUGaIrdS
TN0SmmWMOi3VDSJRC3TjBmWfwg22zyZBX7fYhKornWsTtVxxoHpsa8ng90VU0zIJZXRCn/0fbpVy
eo/FExOZ0jvU7Cnrp8UUaFXX5FkSdeyE9rgo5Ef6KTHTCw52fq60LYVsVzFT/Oq+RnsSrp6D5hDG
zwMlGvV8+IJno+btI8voiu67d0ffvHvHpqJCQKqFEZzKyofbXN2jrtJ4d/0quEhTOMgVuQXeY9Gv
+xtNNKIkIcWPSL0gWrOd7G/JlWLBi7eryn8w4U+0tovAqFt18U6jQQD+Y+wIjJeN5BKViIZTdY27
RXOHcUtg8Lv6RQXkyK6U01FEnAPdnlrYbxTPptzpAV4L6KRsM5eKQRBe97yXBu3T3vycYGQtGfT5
ybT+Aba5pBfhuDRMfD3ZbDIBwAav88XZpeajW0QdSW9fLdQRsLU7yYmOk5HaVEY8bnwJzqqzoGud
+J5OnD7W5x8zYQzExCC1TouwPR3FvQTQF+u4eW9cGSWAdkFCHeQkn431Yh1LDvgBVytgyo7x41aA
iU5+Fh27yksrzECoXmdfOwvIxeoXGZ8c/Ft4pe64cFx0i4V+T/E7JbXqwgDAbWGLNKXsCZw5XnLF
Y5SGtLmaYAMHkwtyHfXvGQaSqH7w6HxH/rsUOH5DhSZGPoKWiiBVfy8GGHpxvWClrDcAcUBZJ7WR
lPWJhNT63+7xFYJOQojV3q70IKUEVLXoJoJ2LPe2xQZb5acfvlAYkdvrZu8b/2yUCXyN6wtTfoCT
KAF0jsAMlbeeuFzXhNLgbd7rF8hD1G/PnszyvqK7DoRYYHUOpa8dAzp5GaJubG89V2RW5rR/6Aj2
WR6BrQne6mC2J+L2Iv8DQuG8Sdl+gXyU1CA2JPfaxu3XeQ1FDtrFu3WIl4pWCc+E2Ag3smEF3Ymc
W6HXhCP8OOQ03EyAaHvQzpdxkWBqNc+8mtTuMBlimdJFc5WnwhpXt37kTI7wlr4eBra8F5n+qf04
Cp5asbjHR6bMeBYAL1UyrIARPI8mUG8rUqK/FCllY4CkWG6MYPeHf1KzJ0EcfnH2eBePPzsGGQ6A
BORf8e/SqvSzETs3NhxKdJqt0kcrDq5QWiXKQjncIWY+YywoODixalRE9X2LzMxf7kktsIzWd+Il
4aqfJadNuNcojVT7P4VlcjG5hB6j5MyyzgircOVHbTn8W+TF1X1srpoCDiLQBabhXw/FjMDkifF9
b73GxqM0JoVstaDAQbXEcoZjmKKdthyly0F6ANcTCoKo2C8hDTXEeGQWZjWs5bD0HbRppu8Pdckh
zU7ZkvqoT/oTjmDnRbRkFIIVcmSZqOV0CWC6BlBR5NJuEFQ4dXiNil5gONVDmY5hy8ifdzS9nGTW
rxNJBKmmDSecUwOSmckp6ocK6LD1Mx3BmkrS1mjOkYpo7Z3nheg1SXPYeXi1DN/G7lK0GlsR7TCz
Zky3ZiCJDQcMRJE9IR7VWZe8SG7SwEVaGt1EdXdHi70f1o7U+H0AidSTlow5LIbbQaRhOJrFZVVj
TsTl9JHxkFa8LN+r0LHrx4FYZOT3l74zoWdD0Al5/ZL6xb297xgsvAIIPu35gzOHqD+NJm3LIQUF
NrkT+HEzUtCFaQulQf1XPKelV1BGE9FXYR6Rqxgl/NQ4XhWpSGCW61n5EV3NtU1tsa20UpVYeMtK
KKEwXoulncbLWjEytLP3qf4qpEd5ZbTdbngu2fJmT1NWJy1kPOKrpNuKqEqYj6Xq+LU6cgRooj3P
Q3psEGeb49+kNaX+J55YiETwx+4lDJ456FfzntPh81eAdS3JnuLJi2btf2MT1eK+oFbmv3+rTn11
cD/sejp/zgSwbLiS5mjC7ooMxiyM1PuisBN1znEX/agSQ7Njg7kQd+SRF1RgBAxXm5ESq4wBn2gI
Clz3CV+w0umnO6r/yjna6YmHLb1NcxyZKwlnKMDNg5rEacxoCEJupt9f11J7I0ytTy3DKcdNJnSK
AQ1/OQtypnGarg+K4QDnDh4YHUar6jeA4Ek+jnX4MJC9ki1ULgAyDv4pnztVo7flD3ROLPRUdtOl
umQCQz6TCVOIThLfdoWMfFasgqK9wz/hfM9yEsG8tiJxJ11q8K3RrfcAMgcTI3cM6XOz8DS39cJR
NbwjPk/773h948W8cPaZ2SGoI+uRh91lYlgxJe0YCrhWk1vwusBjwX/Kx8ctcvNT68tF7zAd5cx3
yeHgpeuEwcfyGoSZieTKMv/yrYJI+Vxvz/+uHExVS2MQJRG/AsAQHFforbKXwZL2IdS1j/XiLKLI
8kFdpsUU1gWCzSuNLpOhTmsHcVo/MnJlH3w7lz1JaXKwBpDoQVir8BP2rZElFPzoCrcYfds+8mme
YVDyqYTvLUCIkTlLILZ44YQkEx4QIRe9jXjSr5+Zef9Q7NpYYSvpfq6YAcQw2+OylJFozIsu+CC0
5Y8GXcA0+/fKpZI7GrTu64vsf91XQwysnG8TdJV1UYOhTzr2uVR37SfAXfmrEHk6AfSRBYRkk5mk
yvTrOVKn0Ciewf5fxj+bxnw1iklOipNxhVIGY5OnJUoBVf5qyD1+o+v6RM4KAGpEjhRrSHbHkSNb
01bNesEL9ypZCA7w1TouW4/uLKpyAno3LhhD8GNpaVzCINBsOXvEsf9ed7v7dAkOUra9IzGCLv4Y
q2WMS4pPHlAztwEvMGzD417XO3Qqqq2mBFzsnlPlrje1sy6pqrRRMDdsCe7trF+NlA7ZfzdW/i4B
3HbUSFl5Ky+3PYNPgolGmSZlbZiEoEl8Ed1tB0V7WEb2BOavQqKnIV0FHkACg2HNn3MsTtFmAn2A
cZiYVKwucA6BAG2HT7oh92f9cM2lCwqKr2t0vbkyfztT8QsXAZr1pXhVTA95XYN0KjD1hFqSeoeT
taRdEDQIe2Hiya91On1hKywNd7ATgRDPK+op4NwLthqxugr9hXBjtnAnV0RDkVpwts37QwWzyVQz
q9aaPZyWp6lGsZFYO+8PFibdHrorNpRMKnrMuHE9YotQNxFQTpnK8qhg734BkPdT6ZEyv0txGazm
RfRNwsE4k43ng2/eVTVr6xVAQltxGiezNB0Kwze3aUPU2tlPXFOt3CC4AQhzMhsASUBdB9KgMcyW
868LPgOPMTGx7JxNUnLjD+7yV1OCQM55W0evsb7PXFZ1b74vqwB8ZP86wabhf5F+qM9fyfkeZ+Zq
k0t5RHWonBV0g9rHfuethR0+ywLqzTMjhBWK7b4VixVFUvmLL8qeTbWCeyb4gA0cJSh+zgu632il
xBY4suV40OPS4x5XTAep4IfxK6uWHpRUP0f5IiytXpklq19cP2Vh+RLTc75m7Ce1y9Zge37VSbuF
QYlUccIXZbvwCUpUdfo2hgnHQJmdQ6HnskHblxefI44WhPTmuopfcDYIgJUM2B0zNCXe7ITtJEzk
FrEW534NstHKY1MV+tlwQpK00rKOTaN5EpEeX47Gf7uajnlZZhjUpMGhfDmPsFsosoNyDnvVCGlM
p1qVe8NPyFdF366vGQSXPLM8F4q7D52/tmruvpo8OBekObew0tdfT6tGqM33WR+V2li7MoEgXfJv
mGRYiGPAGU5oT08yOLFnzB6rWB9DHCKFM8wvQ3HsXpBKMpo6vSDpuNSL+dB2uI3IK1PpszuxyKk3
augxXCAOLSrjENM08eoa034wG+8EZ5KK5oayS+QYBorLFxsnSZve27Vg5yNMQA9GIjRnDxWOYxRv
hqylaULwd78yYcJ0vXovdLF0spOf22XFezj3Lm5Nlacwnpwdm7yq7vlLUw4PbQFG01XafOC1ywsn
8h8Jagr7yRF9COx5Ny4gIAQAxGP9sC8CPAnn8AI4ipA+BLDPLMQNY1295pdvMEDW/Ck14v3ali4l
AbtJc6T2mSRXL72d9koOG5IHE4iudXFlwMnWWm3zyQN/j2kdTaf4SXBQwlQoULgn4su6Gd2Jw4nt
hpnbgjoAqa9B0NENrjf02xQq4VR8HmbASizP99mswhOk4O6RcQqCEO636iCVZ6dhjkjZax+YMeH6
32A94aeRmSUi21LMGsf0sYTQcwdY21tlaWGUf06yaRSCxMRFpg01QeqXHPkT628lNjUqgXnRqYSJ
xn2qdWf9ctcsLzbu/kTt8/qvdsf7taZmUxo+UUG5h/qKMVHJ09hxq2sZ5N54o3kGGiIN1RIf/gQX
KY2QpUuDQeeXe/343TPtqzUEZFmevNQ+RC5fZNWpGP47MK0sVXMf6s5ZMF04RLYjGMRlKJAOI4nG
rq6d9k6JkBvQl2rGgibDGXadF7FiVNbqcl8uL22oS4pggQQh3lZkRnuAGPh1Cin0zlW5pkbSLK/4
UvkmKwNTz28a3fdd1XAQP761V0UHHEVBnvJjDtKxDxHMVDBO1LKVqUbXIkSMFuQIfs4XcrNjslUp
/FuJ1W/uNlOnrihEAIClncJK3yk4+SM6VJ1r3kdhBMe2HZrd/U1NG+4z0jdUETMtbb3FexnkhT5m
AOMY78rDExApQpTlS1agPtEABaYYdv1drL5cVkg4Vw3IajP4SSos9HA4YEvKyx+B4mf9C5WsILmK
wDUHmNfbp2fNF3z2PtGA1Nq4czw+QN3hyLIMfK0OE74YcUKF0uQCt3Fxz2EVb2bJL8FrzBrg15P4
qckoNWTqpiBOlrgW05Vusm8RAfSJiE250GtTFZkUE1KSnDjFgQcnnpv+FS3Se77wpr7okaDMN0Al
CpxApfGO04Gc9kMXeVHYINwZcIFOl4zUwJFYL1VDvdzUqLTCno26uPt2FA1010nyaPPgxOJuzAHy
LxPPiFRjQatwNA3iMpTe9/OiTeeFD16daOG0wpKhqmUTil4OCLxnBCN7zxp7ovj/nZbSD03ydpUS
vEZVTwchjZmS3m/1v5daz84cXVv4vhaXqMzNOvaRELGgzpzAkhbs1UfBEgn70R40KjKawvEuyEKm
unzB7l1bdINJ+pbIlEpFcMM1zmb6KbZGFt4GPYlIGxvZ6AI6NKXEQMKF1B0X8RuQqVCIfr9aGy/g
B+Dyr36FAAfrbhgAbExR34W7dXvKJmpsts+pcsB7wiXX6paBSU5Cf6z2MoK2UmksAGD9tu2+wKZg
7FGUwoiASkm0lKBGBUfQbuQ475hxjzBxZeqmjfHEYChscHMlJS94MW0WUPY9UaEZaMslBYP52KQ7
7jiZRyshcYQaNvB2ieGXpNpXvRmhoj8EHmeRfezc3y7fabUBb80iF1ngtVlR4AuT3Z1Jx61qNeVN
JfmkApw+QZhSmqjDD48JVpZC4C26fYMfDdAj9SfO2MKS9g+3OsHZqXOsg+MVlIlncrm5uy/gP9V3
pMA2FeyTW2PJNHrZSvVp+UU98vrTPcrvq69llQW0FgEs67T8Yx8cecUwOuyFJE3wQdCf17P25EwL
GppTa1fGveiZfEmcUkHKMHclRe0S6Step/KITSnyK+OB3IBGNjJ2d/Kes/FKTpZ4NLubFOw7fEMY
TUmBr9JywIgERIA5aCAKmSAo5g0eAD+VcTgvGgH0QfWB7JlAUux6VoJzYDaM2I895sYmo/OAN5mu
YDNbSwo6PConRnk3kIjDBs+lRBTIn5n9ixGA+KX07k7xWJexMsF9oGqhymxWZvannjklIcG74Jir
Qk8uDZzB9A6wVneLorMb/7EN85o9c5E+gC2U7/kVAZa2uiR/BcjDATF9emubzWCimNV+n+oJ0fCr
8D/fvnwn4agKzfxBo4JRYh8sISpjAbuAUfa7sxgGGrO6VysDI0DKreOwFxZATn7OUSFWs85cAsHg
NpwKNUttCSFiJYkn8Ha5h5t5tQg+Akql8NZ7rbcA+PYi5A/QeLVAM1zIG42CTVl293sP7+EmkJ0h
v3zeWacswZ5WVpP1gOpo+wEBryzChp8wQBBPdXDQwzZHUebcVECFWQNqIt0HPekgqfRr+NT6XQ4h
rJmvYKDSBPn3BHgvvqWw2TwIAqerAhoqtpu9ZBlydJRFBVVmqXkcYCwknHzMln4CH7q3gDbVlZ7O
P7IgGpRIZw6TKWOqfmpcN/61f4w/H25SDVhlC03fV2eMLBxJLuweHBQzJUoXqzEdOXXoXdwgMo6j
8f9RAywvAVC0uGIhsctLkRckSFoCF0FWrh59qvrB3cQj7hJiG+14quHJjv3sTE/Gt0+/YZVcnK1S
hEr+ZMS1d2DNP9RUeY6JlM3BHdZIKrxYrtaDAi8E2aNWue5Py6nuqQmINkr37BYiKw0XZuqjxZ8F
TZe3uhGdvUdTP0y3LH6q1hL/X/rMVquMwymgYMfmhpYuT4TG7T8Dlvo8mGC88bre1D27962H3Ukz
rQ0U3e691O+aqqUXH/CDFzC6ZLqY90UA8judfeX1KStqeZf591kxJ7Ab57DDBdPFx/HyCybz/af4
fb/PETlKj27t4L2e2pXST/m18vcLV4yDrkQAj8tH/Ss4TeSwX25tA7cvtuN4FLRwhuMbPMc46AFq
Zj9WgWIi0JbroSteT22+nN44YfxvhM3nwVmSy1CuA8qU9x2ByfmcRD87bGmRRfkWGPw1ukF2J7uN
HEMve2Tpgrqi7w0dOpEw3kKjG4PV95TO+foi9MZMkH3e7xrCCkqqenKReGlOl+LPgQXZ6+pLbVDf
Xvh34s4a96MD2gw25R7iBnVVO7auMbusht0CTlEoKHzR5NiFwsKyGou4znz0qwr39K7Ekre1SQlf
F6XWr0LhNnpkgXvoTYCZVBOJnt+/oUDRqBlfDirXvH+90U782eXWAgTvE4eVQHSU5Aj3IQfkkyHv
PGIwi46zKnAwKzr3nRjp74J08cWwiuPPqd+6DdP6EhOBSr0Cftl/Te3OAesqO18RoXlx9AvNAQ6G
ntd3gUdVu4a0RL2xpyvL3VPyU9jecO+KaNwpWEHPWg9Rl0J1RpcgdNMzPevuC1yxc+t1PIBq04mj
rLMw9ph4XnDk0VkxHm8YdHBs5R9NLX+DQKqLpXxFqXlQM5Z0eVnnhge8oAl64l2yFnfONBEZqCJN
0wK7zqr7f1AXXrE7V8AyzaE30604D2v0U31ifdSJMAXfbuq05XnxPXFT+Fx1uU1tP6o6U3S58mh4
ZIsSASAwZrmOlnRP+8z2slvFemHk8/CfR7miE5vu40zsaNBq0RxOqOO9mZkyPCo4fCwgulFA9YtV
dSk13Hfc1BAUmq5fnxIs0YQAbuXjuZtPkCn5ay2wuZCxU5aD4ZSRPW3T3DHY+Z0BLTRQkOpFPwZq
+5HDvC0qlwSCIOvAojY1eVw/zYvcRDCh3uOc0VY8x2r7wiRS4T6hjucmjQEusybWUfLd8RoKKvEX
vq662RyxYYFIzLaK/yfTCaneJsscrbkKfl6ASNN/FD0tcqmK4Sv3s6Toygx5JMjsiU7ycoH8/lOi
lh5O0bXYluHlJxaCaDVAaBmwDoAk+zMEBVwrGNG6diC15NXj323COzB51hBk1+y9c+GV2KkeAhSt
pi4yTgkfUqtmMssKeMn96kLgLg0cDbzuuwpOT/gnwXCtD+TxiXI7oI+rsuyfEgshF9HzH58m4Vg6
SDXq/EQwQkX4yFjHr+yyvFBYE3EnQGngjvbO2w1pHZaKzevaSRFyiIKbAUM7nJxDbGRVV/qCs8Cc
pCrE2+VLZCdMBfjXgMIo5/m437Qyyph/bcMjWBzofVKqKM8vR9m6ptM7AHlcQAz2nJOHreg2UbUf
rx/Wpz4LpygnfUz50W51PyzfDK1r0qclummjueK2wh1/xxgSNFFzYwSa1ps6KNfrfNjV/zTmXHTw
OoZwyteXkVNTceHu8Hfq6z4UT72JDslosIx3iNiDMkKjYhJK8dhp6tJbz2J30lavrjQcMcsq4Z8r
gz141Lo6AWgCEs3WgI3pOzmoRD7bRHChXmOPkJJnWrWGY4eg6/Y6MW3NLwL48vv5gvkrV+/QXgCE
AedEH+iqsvx86jvmAIHoazSLPEy0QpZOB6SXi6ef3MXYtRPWnZqxC7fps19yfLnQsy7MO+p5ehpu
r4MGAc1ZgGteNL5mQANXFwn7RZ3RxqkTzXZKA/bzWrFfF6UlNMWsRavnI6ZNVxIBZWtETVF0+Nza
MWzhZjVp1583afnuYDzsleMi9VUjHeRoNmbT2MUhoeNA/x9gihQhcYRPPA6v04Dy+GdXadq4EpCC
YS3EmyHClsludjZMAulWWp+bpoiLUjK2K7xiwH6q0JbOvTBxt53VCSusS49tcaT5/+tn+s5fG6IM
DWA5Q+j0BTUBrhm7qNssIIYG0zRdotFSmYkR1dIJ2I169OnvKqGoyZosTLtbWIEI++LNdvfjXGH4
cf9PtQRMRj3eg4t17ltFY6yNKQArsY+BGy+ElZtiDtu6zkyI21io87Nx+sL14gI3537pfiDlCT1w
ex0cT/GFO/Q4h3oS2rydK3xThguzmHSMMKVLrrxtKcvQ8PyVoZqa8JmVHbOfKk1tGndtJttDrq/m
LGP9/7fej200Vkw3VBJuusPhFEzMJqp5FVmNfXikJ8uqL65i7JGuXdYM17aP+/xjMGUowFvzgijp
7ASD6fnnFuQTZ304fbaoVqggQuYozZisddJvFlrLTDZAJE/5KHVXVexkhnKKjUZhoZJSG6XTfTPS
P1ixQ6aA2lpIXExvEQ2Y8vewctyjQCHy7rB7d4hCf10uW8uYfthcIixrnZVeeytUJCAc3q0t6cGG
nPxA5BQWUA5I9PvnjHIkXXf60hDFB679FY2U70SciDXOdlYZKdDOTp/0eDGq5z4AZz/H9lDR5pM/
75mM4bP4nZizQq1q/9Or0OcYJz7MVjQIdM67qGIjjODo0fW8u8wc4L6wfhO6IYDBSDZGew6kBUw0
jB8lII6CFVAmbYMOH8WRcPyfF7R9ytADNTQLn2qm3YayKNchgEJzBmDykgGZicqPVVFg/+qp/OIF
sVy5qeVQ9tt2lze+DfTCnBp8CMLi49PXj0E0PRyb+GDHbk1lIfarf9Tz30JqxevegRMP5R0pSeqN
IAl8l5pC0Y09bD+X5r+pWGVQJopG3aRJKrlaGQHDR5aAZFR/R0SCly4PlYFUMIy8M3p0TfD1P+4a
zKIfbF+d9ACXZIfG16WoiizB8vhrrvO8hCReeNn9ImeXv58hjc3CvYBUko8Fdum1uCEls7f2n66v
qQK1Rdw5OtsU1xj9Scg7znybs5nOy+W3tNEX+q8dV+R+DG3VFApqpwTjcDq29Z6KaJ7P6GTJKYqM
U44w1F8AdoGNBI2zux2bhM5Fzqvtn/+VZNefD4MWkirRXJRHLZAGXVqEP03UXaGIh4M19pB14x7s
+3j6oVpEcsNQqfyFn7dFFNgpUTTsXEGXum+vad0+5vFdPcdA4PJ5jHLJBObAMIjwuxjIsAQboc4B
/8Kz3MXKBUIjJQKR0X49AfwWebDlKeQaWIkoze8RZAVtHhW7EaHlBsbpsS7Il+ix32j1wJbCMIp+
wKy/uODf59vQ+ksMGgFcA9JiMMqilHk3kd3cco7Gg3zuQSehcDza/M+F/FnWoqXyKo2dSBrx+zbg
kXlhZfcmBoc4U57ymR6cfL8a6gICc/+n1+d0HPlM9WnfD0tYb3B5l2CcjfTzc4/jegNGq7G7noK2
WVvSRpZfmJw7GE4zou/pUS37HelvP6+M8u/IsqWWrOnJxXFZZh16vjqldMNoWFvdQImChnbK8Ept
86EYIycWsecEnCaQgUiTDtLrXaWDCGetMO/Nqkn1+K5V9yzsqlxSttpVeTKiRWTXdeqDDHh9wo8H
Wq60EpKsNIfKEgiKEw1jbl37HX2gZ2R6knt5fhjPc6YuNxAqbZW5tzeWleHRgrSgMPWt+jHNjH2w
YxoTU1r/mqs+R91mNls9CkiythAYIf/vQop67U5Y8GcxV2mVfcqnPoHyz6+frhi50XbiQwlux6r3
dMxVmEsqR98W63OqX0k1/uiHoe+orbDPIuuD2na9TCHxUSGmnZNpU60hW1shZOjCUG01oiO3kcz2
To6z3SENDkQ0dbkfwSbsdQ+2HFwU/8pnq1AZj7lF7qOM8x8KwJrW433XcOnWlVSTidzGraXEpOjo
AeCHpx/3fL9Bbz1nt9q+8h+cCE1qctsmsIiwSWao1kDYNa1XQOnQ8ZvaduSUvAsA8AKQVlC3FVH1
PebPuFY3WK00k9uJAMK5280B56zoQkIeip31lOakAGm/17JJ7aWY6H6FwAE8kL+gx2Vq1y8whtiA
qwwVAgIXUwf4H7elFmjfC8SY8LgJNzmbDCxcOidM9PC7cKx4QMg3VXqz3/a+TMqexrCNHZI6W2X3
rMhdYIK/8UeAKnwluR/7KmSKNAVdhEvnyvwRrI3qDr/GGBCW78zJd4t3NPzlqKJ7PKpKMHHs7oLx
J9186tYe6DFxiQg/32cpvONHjoDKz80y5yUhGzyaRVDVZa8W3itRpS1/eamyR7T/eervgwNDnj+m
9vLqr1nX8zv+3iXX/GqXrYl7SC5I6l+JjRo5yK2nfM0bb+hAQyDdw1+MEZ7saldyS1TtofI8M0pW
UBGy8qfc/Nx6kR8UehGSZGQwYmJqwS9oRrAlsnuSyTRgwaSsTOOMDbjHDOWXjudb3Z9Jcu4B2Twt
XtdbhQU7DIIXzjeYfcdD/dvfMXisBOdLl1vBmav73uHjEDpATvmIKIjiOgpxmvS3vc9WZ9N7Jb8Y
E/lVjbIfZKGkQFjDYCGyyRq4L31Cze4ALt4lTPFXXfRrBWGEVZkrS04DIU4AVn9vr1cN83pd11fk
7p7cWVWq7zdimmNxLsB3ZBmFvwBiCl5Ojys+DIgj6UPjYkoJZkpXNK2UJ2m2xiwtsxwsFwqN9Gl3
Xy+TtTH/7un0tzN74w5ItyWCU6wKJBJXN1cin+zuzVIg4Hn8B1WPrszw/SvZYkXJj2WeIKEwAfmd
ptbwHJkMjrO2pmzb3D0TeknvJLXZzWunTYAKF4fRqJJCxI2oeoV65Xz/G7yjHVuTKpAkHNnPluKB
mJO1ltNuPIVbpx5CBGRvTFwYSUYRQNo7NW5cpeTZBpa+lLGAsDym5UUGCRGTFrRvO2tswGLUpaeL
lZ/rvDHKCXGwGh6vNrxtP3o6frTuNegD0c/fN8BrgwTZnVfSWySZddDDIxfEGteeubR1z1eMdlol
4CZ49AbPzk6FcoCIHr3WqVEOSgvLTvQ3Niicwy4ZHoJQ10XXc+09EAoOUzXnLc0vKRAajA0g92yj
femx6+c+hJ7MiBaZETkNm2+iYfxSJDqUAFV1tS7zne2oc+GByvvBwu7mtMHhnD09+iWZxXMRqZNY
A9wtE+L58hFcXLmF+P36ETweZbcbFOrtYrrQDkIhft5EYc14iG+6N+xuTeE7ss3ZTygKfRilXmUS
jo8JmXixu2By2kkKRNfe4p7Vqwvd71/nws+9RKMllWS9d19wW5J4sjfLIJGjoRWqMul5nppao6G9
YaKNzdXUrQNM/TDyeQ4sm/Ri/CGcq8I6pPPaiVp7zaNMlPVcHE8FuJiHawxZvsdvfl53nu6qBgJd
Z/O9/ZimGP0r5/MVn5pSZKI9HOf81b5Y9v78pMYHA/ObKSQH+qQ+wq1f1EXz23a8NoSLw5CL75VE
KeHiVOqC87QwMeRqghfyDFEK/b5vZyG80mgU8RLJGFMcbluSS0Kvgoss80aaXpcxzhYQ8e1iLXYq
R5X4PNIdOXvrnHZXW8HAxWavxXm2YJpoXmvTw7Uzr2g+VPuQGJHhQEQfuxz5kgKx/81BKPylSP8u
H/ECM20pMo2BKPwBLKc5opNQfDZQj/sV+tTY48PEQzBwtUciI0RgeBZTNxGI0KEuQ0abNSJ9AkMi
pgLtt70571eFT/soTZXdvjWSCkrCroViAjjx6rfYdJT625DMvxoKE5bL69yMVMupx+Ro7Lr88Gs2
LXWAfGiaU8QPrIUFzksonMLWyWx7tUYeCLDecxpTEu/PWGDvjpRppmPdIha4jXqvQocnejr1tk8B
KWj8FXhCC7Fibswcx32oMCrKAGOWzNOq3QD+rc/N9odwyF/EtZ2QrzTsV2CLmNXnhJ0UU9kAdpLk
RFgwDKL5TXIrOElObANZcPt36q/OVIVMxmYulZQ3sxKowbh6adPFO/+1BBaX3B81cLQyQtB2Pr9V
b/CD+GbK1aQo9t6pPayyCqXx0xnmmAE0xoqMvZmcS5lwB7ogSUJTxmWEIX8kdhGsk2BF7sy/LIYM
sH/srdOp1u7CL1zZR5c6QX6TYrcovrXgXbQpqbghuuVYkNufq19NlUfTgTAn7LTN0kL5L/U+tCtH
UAxx1gwwTIb2HWeQLU905ckncXntZfelboViyflRRSzl3ODqvkJcdx65HhNDSFz4wFHl61/ntXws
MvyX3Zs2m23HNXSgmxaydrxFV+I/vJ9hPgsL9pvDYFKz6Va/WHw2wFgPCX70wl/7bSyM/3zsHeiG
ugCM4t2YL/zh6VKH19CntNX89ZtkZT/1plxPFvlPx9toHNIbLLpBmDPjHiowHApKEGQ4x69tPYKT
HMxA1j2ms1K/4avr1Fi9LVPXFW2jUxIZgUs3LaVM0HZLiPrDGyNgW47YAnm7FfrnZTjivMP5sWs+
b74eizpWmMtU69f/95q+1o3gLXd3Z4O642wAZ6FptGDbE2OowfNberjwe6k8Fvqlh0Ks7lCo9wEN
ShtnoCe69BNbjhJKdz3cNvK/45dvrrFSs1Lih3YRi0I5R1Fj3B6btyGL4NFPWurvPx/0o8Yznuc2
TyeycN4Pr0/iIxHSjnBX5fLFtBkdc+JYFvZcb1dkLYgDs2CSp5vdvSUPH1kiear24NQmZYbmfkVv
xnrrTFE/RtB5PUZ2lbLNORI8kB64egPAZRT4VCjlNS0gIS11uyM22V/xXB459I/xBQXXN2XEAosX
n+aKZEQ+w2eA5IeAtY4HauUkgMVSRNXYuIyL6XxXW+pOkLSSMV/ykzAOclJVjkTwz/JiPEuT7jzz
21diPE2BBemoP9W7/2B8XICN8wMiKWyRmv9G1QJYx6or59d/uELtSt61RNpfILK8VY6ZuudZdmv/
Z0gsL8Hhc9R3ULm+Do0+T1xyVuavVDgYoaooawFlVxsjj7Fu/B/o7PckGK1vYr0pD0RgScW4sbjH
DgXUyqQquC4MnINK79uaABc4/ZpsOPuHRAup7Y/Dib1Ced5zDV0BMUDOjCfESv0h7znqL4rZjG6W
q8uN0CDz8nlCDt7hXGtDEs2WJVmkOx6PTvEaxLOvRbcqvou2Oo+SLEUdc68L1XMfFxjFa9ju99yP
2YuYX4Of01rV9bbwKyzGE3xPQcSfClToicKC+WtjPMqyxFsS8feOk4Sm/V+15XtjehdPSBrP7mMf
IwEQycJ9PEXG72/0yy6ZO/l+Lt0JdKB2AUK9ccgdFAE1N3LGiv77BAKtf/jLcBjxP4eJKMDRjr3t
fppWaUIdop01zUl2TciqT7hVQMZCcRK++8Q+XVjlgntF6+CHaPABrfU9NVHTNsZ42BQ5E8apcqzc
w1nnGL3iLG2hIuBXW5F7xa0ETeMqi9hb9DyzlIC/8BtMN5V5wEHiFe9CTW5TRjX6BkXsNzDuJud2
5FJFm7rzC18YbRRMeoKzGR9wLGOxhxZ00BSkZmpSo1n2FmVvJcvY4uVa7Tt7E3jm+KRs4Xr9skXN
k6OxF2hdAQU2KyHUhKKJRgEtVTCCEGb3fzI9XlmbTqkXXMNK5hHb5AEk+ksurni1f0IZEnQjXtxF
PPW39XNyOOSfrqZg2odeCZtv4Kn07NcVHh/WefZAfBfLyILqPD9UnD7t9AYIlj3d9bo3tjQp8GAP
ZyJ6vPgJVrLZ+uF/CZifkFRU/jDX/Imsft2I4Chbn/fK7OKF/rbMsgXA3Wek6uwL/GWdzZEUYNuZ
bvbo/dLHWzZ3Rh5F6FSmJE0sgW8zG/HNFxcMVbLsTnDb7/7WH18geWt8nEBEzvWJjTaSuaAYd7y5
nxANoyx87/lExBJxJBwXk/xd/lUmv33dfSZK9gAPrGlelutEd4R9YxzW/jCy5tkKr9RVohjR/RB/
InNYNt2NjRuPeDx0sc3HigromQRWkE5J71cuVx5DYpIC/WkRB1MpmTyTSzqOnHP+tujzOXkKVIB8
iaYxFyeb8G4rOgcj4Y9734XzenmcVqn4zGpt3xlCnyU86+8/bW9goiouX/5dmYpt3UB8PkyJycNj
Ke2uWNktVHK2m9O6QhJXauLJt3mPSAQqsm6rUSPeG2IvgB6/iNwx7qcgWm3xfz+N77IVl4sOGPIb
UeWqgIyI5t6Zet+Hf1fZpGXpxnm1aLFSAP+pDPzoc1/SksQsmzpLmqK4Jc0xqic7R2G9DoIOzI2y
5MBMj+Iz9zp96IW2wdpPS4n80abN5tRyItH8O8qlo3WJucZSh06dvURLtVpnJO1H2HFphAom9/yy
kqlQ/Ly5uPFCciXFuNv+qD025tbb06Hp9i2J2oscR8+pL4dBt54ja1hwR+C6rg4+779GO1ok+rgw
ihobe6/wq1B5STlCXHXmakCHs4i33j6TK37Uz0HKp5LF3ozWPw9TthbpFpdKEE8umqY7FIGwjpjn
4bgj5wnIWr0JnVeGt8K2q7AZ0qmoOSZZZcpOkexjWCcx+8B3xxyC4kp44ODYdGrZMmULXEL4v3en
Vs9oHS2XehYNxwHahB2aaJFzVFwddxryWOQ4Q+bbJvYCwMW894Tq59hxO1PkXXPq8esF/CXuAkPi
dfgB9Ya0yl6nahp0NtDef7xJMH85+fyNuI4o3xs7nWCc8hNV4JF6i0d/KPeos0JNiOB13BjnMdBm
3tr9GjqX5NCkdPkla9perACXqI60GHfQW8NwGzDy09AB9XpMMh9f5VleBmctw7fJclyaTONIxg81
ulXns1qpwuIaSjC4dHt+zey6uU+MGodMhhxoYIBY6GQg/hMZulYsW3NC7YNjzpu5iKsEjxIVwdHP
0FbpBXfqLOPgaZIQr/7vS3At8RT4IgZQ/+977djs4gNVMttvzNbTasSBnec1b6BZKuOKTVc0yHwz
pedgs1tDGnrU4xTWzQBajPiyiDKY13TgPzVAG9yKztAaW/3ry87Gp/e65F2ZVa/4UYzF0QbZzCRU
Qxm07T+OYTUbD5Ztz6yOiItel9/pCIQCTmD31jf1I+gkV4WVKq0HyW40tJef+lSSJvjRxhbUWVF1
9e3aHPfQGp6G0JNZbz5o/fvFR+pxruNq3Dt3GzsezL4g655dLQdLvjviYqwxOPinGxSyFFHdtynB
6uDwvHuygWYow1Ha65yk4VCAU4Ce4h/X8stLYbTjlVod8spDilvmF+ogge3WBI+58bQiuRQmNzOE
7PVxJGW5/U+OkmlFErW5UAUqlvsWOPOLx3zcCyAQee0ukpLMWPL6G7PTxvKeRQtIIf4hpCUTvnHd
xdMCs6iuHDVtuH/w2nuFPOOeLRPNO8t0smH88+1eJcbsGvtymavfPkAt6Ppn8QEsa/TplOQeZoNe
c4AcriFC/AbZ6YwTJ96E33uSB1b4z3tUpIKsVHee/muEicdsY5BRjIga5MxsdjamxHKRITEAfseC
qY2Iju5Raf+Ajxr4EWILuxSCWspl4pNUn1TA7WmCbM9GwNu0E2Uai/mspalhQ9Kltx31HgS2E1Hs
wR346Gj/gJnXvfkuzDqLM/TY+n82sFocmY1RdB+AY1l4wnGcpLMCkEqued2omA0dl2da48hZoV51
B3Vk5HE3IzXfENPlsRIx7fa1D+NKIT+FzISK0M0Xw7RN6PAT77yipwX7FYxtSBFSJoap7IZuTTMi
UkQtvq2c8vQUsWJntDJsD6sx/3iSwW0xuHosBnbIiLD7KPDTGaT39SPuI+Xj00/Y7/8Y/mFj/k6J
aYhpt8uKXohsY5RKKbyAqsDSiZiXrQVL/5vSiUaCuWxEEpm5BphME0xB8nqzH8m41ryrM/kHxmJR
8RsVK4lOvEvqrHOS8BDL6iOB5iDfz9F0DxwB04shNIxswNtIU/8Qls92VjXv68N9mLkuZ2FBrXfb
QNVzu41q05NeVFbuOdejx3C7CYRAN45DQj2ZiMyPFaSH4SeI55V1RFLnQg/7kCpWXh98cyvG0tgL
qHdwodSCPtL3kBIFbdsxi0KA/zQtS90hgveomwNGLRDdWnGL6OMwEI59BTROJbHVG2aJCJV9Sj1i
zeS/hzGKQEqBJ9nMu8wgQ48qlptjjYYDhb+pb2KpQOFhKel3JqpUe9Dwc1HARGhwTevt7Q9F4vDR
3r4sMxkeBfE+Nyf0hSTiVpUaJqxqKrK19XEuEZKxAiw1GwX0SgQFw+iuocAF5sKydas1iWsVtbDt
9sxr27wpTj9IiMwtoqlMVrHJ/1t6QuETiFvBPqLDbfecV9LQqzW9arxC468TuU+9ihWgMPkHxle/
kO0rTyguZO9GW2OL6LymBbffPVgOraYFfkb3aLifIgFENF3Ug04iUUGwFoBo5rSQxaYEyslEd8yH
gL9ysghv9DNR/QOt39nYmHw4Lab43cbOEkZ0qUyRkWnKQlRlEtqRAa8qK52I0T+yPEhI1vfTH5Mp
gG/UajslbeGTSiKL3fZYtqKgKVNykM4pHsVWq5vEfA/+SPgxFFMVw06HyY/uq618cx8kSAy1Qm7V
JVWw3O3Y1EWiQh7JQ+EmOZd0iOu/rBSTLH/VhBOSdjkYdelK4+bs+6pNtP+3Zc6xJPdZyKwT4yyI
pw+jHRIYaz8QL5LCC0xaGP06FSHCRff9oq4lafmA+oOur2Lc37WeUBuP7XTvQNMJUJa4ve9xZl08
jD9nun3xugugZn2FOWD8XSDxJGbkAtT0djIL3AyTCb6q7FErA0RwHj8bLfnzjUVW9g9bMp9V4HRf
OZZjv7cqmy3Vft8NDC/4AJsbwuDmBSU9nZ5eghP8/rADqkxWUtpIYTQG9fUxscDAeUTLt7ct97yl
zSyThySWVx+IGBtyJ/6WHrxSMnCE2145AFEwSFNgMv4/VsYl93I2X8j8b+zuIMjNfGMxRkC4hJV6
PCmsGxNPfpCZYKjr7+99N2c6tiW6klJFFdvInnv0naUrzTpYP3lqD+BM/+7GDa529BeJxRtdqi1C
tnrBIgA320jgEqRunYPwsWbhvTOGsdAhe59CtP055QDhPHRNeKljiXUZJElcaG34l3eEfsL40/Jx
pCSVJ6RWKbTwOJaZyTIDIS0u0JC/u5x3BX+T3gnkpmwyAqgL9qoNcSk1nz2ceII9/6olUSlBYFVK
BjjMlZwSn2mx8G5rfi8HuSNyHPMmmLtffdVKAxOp0nTiqr4hFSL+hkWv1MrNaHxE7n7XjrYiZbBH
f5sp0khVI0enC2uB1yFntbTDdlytE+92tK18BqayC9ETwTjM5RGLCTzv2m/QazdOHjAAn9OqIYhB
9EMjFoUq2X6VIv5HW+hnDcLsG7gvxZRGMtlvXDBwIk6T8jhsesiJv++XOp9TBdahFwalb0S9ZrHw
5deKKKwRQ0x/lDKRUkZLdQTVzefnLj1kKQZfqqHgw7TMrAO0Ng3xNMS8TehZWn4H+5pOdWTSd9kF
KF1aiVI9F27+9snoV4EkuwZtjioUGAkVilrTCEMZUAWrUWM7w00VEr5kVQnWT5+/OJN5eD8BhnCa
JXYt/ELoYK4mdT3dnDIcC0ZRKVhZsFkPZZE2YScpAwMBv6Tpqi4lW+IIiF3+FU/5tUkvHXYzI+Dg
6W8ES+7KUzfwGeb6qxfC/Xh0HCzJj6y0SCCC0Orp8IYMUMLIdjD6nOzgldGgmLYzqyLjY2XsAL9q
XM10swPQKM3h8HVkFD09+WtK4jw2NwleWQZnFih7K7PolFH/3FGCAxBVBZkI4mOqk3XpUrF1/ihZ
t621+bE0SCkUEbrjuxN8JAASvY3hH8EzJT/LcIGw4EhCqkrIdmE1wjRXZhGKyqMpBMhEwSl6zEhx
Hw0HmgtxGxiTbEsTHsojnwcf1XoefHQUM51vo75prbhkXSbChuPAkW3HdZhCEuxbijHjUlRZAu4H
nW7ni/OYAeqeLaLL0pRe2Vq6+kMaGemI/z7d6RqMGYEJhGDAgGfMzbrL78OqkjJj2nFS0jaPrVit
Tp0TKs+6g5xt9GFcJptFUppmdIftH+uWZM07IcMQiEzeK6KU2oA+oIticwCP7DSXuM6/pwXUfK1Y
8qAJGqEX2zk3I+8iQCBAKdFnGR3VjtO39RD1nmRSdpwJrqOFpbLhTrw3Jho7jslyPMYoEPpO9WOE
6yp1yR9X2IYVDZufEGDpxNY7lUIRhlmIV09Sj0F9Ro1kPPGG49ZDrRqOEil8siYh8YipXd2yC+fK
oYS+r/hbQwWL1tfpiKVfiZ1r14dhorr1mwOVwhlodXcW7qcvN717AGIXC9Dj0f2K6rux86VTjy7X
YcfvfXDzze9yw1X2LmSGnNHYASaafe/kSp1xILsmLovqwWxQuZZ5vrIPWCRqlFYweuzKPflsmuoJ
V7SND84tDRje6hfuy2edMjQJ7ykHfxlCWh2Iyujrhwu8Eo2iqzu92s94LwxSLsQ1bS8An1yBhCd6
CFto79qeWHQDyoZOwqltXbQ/uiJuROB7Qo+xMihWbjMu2lZ57ocBkI5o8ojiirKM+gPQ4tByRzge
1VP9pqg6TQ9m0wZhejAv6F0dY/mVQjD819hqK+PRBcK7k7AqdROMtYVth3ZcbyTwlec6MeUaR9nP
s6hzOQHzRElTc2EHQIFhPtCdJ2oLF6VUJRIJ6nN3+Tkn+L58CcCL8xGAJ/47wpPYJtFQSdMlBLmx
rCbcBr2vLJSiU6sZJsQqgnsVxoKZzLRpwllW9wZiTbPC6IxwpT5VKeXmaSlhihIGyCTNObsTdvqw
EMZ1Kj31sgChjVZ05DWMfWq46EQjenDDwtRiRN8HyekDQRWqAIx/Ssh0r0YsOhhJXFWybLlEGUfv
2aluXq7ywpONdjzKsxPgw/VPHdiA7sasDCja0USDW9So7QVv8IeD7JmC5auAloftxL50SjY+W0t9
PgxmKM70zp3BvMEilfPPZC+asIYL3HGj71Etw3h8/O0maRaszAkIiMSKVSRIshdhe4e8I6kcFlRG
gCbU4i3vm71S1SCUActCMifNyNDGHdSF5Grb+ua2nCS9cKlRT4YbBZAQtloT6DCuQnSkU0iK9YD1
XiXRop448wWQ6olitujr/H9MZLnC0ulI8b4hkSNqjDyqFYzCWElFlS7dFoH/IG7I3KchimtYcmI2
VXu+5Dh4pcpGWER+pTFt/B2TGDz+pi3MT+PdSrKSwWAdMh9fGH/WrPnu4gmHshGO0m8ijMP2Ty8p
VLCG3c0fNY/x1VZQeRnSGW73Fa63fXFO1PguM4AtXNKlX30nIV1si3mIgFDRMPBztwplnlh1W6q8
PUN/ZAo6WPdt9DkO+c4s/lhMwxlV2RUxexZitDHnYAE764gPq9h4tRZaRMawGyMyQAS9rG4hWmxW
p6VxxeSAO6nXFPaQO6tPegQpNDX7yrqoRTgaOb0OfD1CfDX8RNfKEK0cuWgQVQfqVLKcpv42VA3y
c6nVHB+3Xn6WZySmVgljzQhRZV5PwldoUp1JE2TRX3hd5BLte0JWdYqRDQrxXAfGTnsS0SPLvC7y
r1UgHOXxFTCPwBn16XxA6/MCbFkGkxiKOJGmYarUrtgYy1g5zcaw7Nc1+MrJJu7GzLePfIReC+WP
0lWAQmtMYmzJSvWFbUEYR+YCrj9JaLyuhSabn5gWucim0mbdRHtevGqV5Jv4Pe0SI/ZjoZRnWY1H
z+CTG8HxGpqt/2dFp/QyOzCDWoyg34jKXcKW1MwyxjnMfsmfXf9gUtGdQvCNFTIUhTia23KRkd2j
bCnBkrkwfX6pNg+3t+8N7SNtwZbFYvxFqZKjo9FTUR817mFrjr84fh9cIZeyr/snTs5RfvukJESd
UdU1YMf+zVVTujXuINMHZn5IVLVDlX9+zAM0U8yqfLuVjBBF65hstBHeI5xw8amSs6bcmuu2dPoH
1EG4ox4QS09R26sWfWeQiyOC38bBP2l9/u+/WDXVWZoTyJQSTHUIXnh0qCZc5OuwR9/vRxhfOvVT
oe++ZzaVdJdXsdOseCYDVP7S64Vr0QBE8x+imwGukJhjh6NzYEC52lvSJNOXwBwJG7Zkq3VP4iz3
Y7P0+EMtwDKwE3CUpftAuCRL+uC6iaUPtjBW9GTcbFLOt/y2nrfbwBJ5bRDUggZf4F64txMb+YAl
GSLtRO+4+2ZnA91Am0K09C/gCR1ZVJHh55kIGkLI25Nixd9hmEb5W0iuULv/QCBgzsHHcwVxtpSu
YWuDwl3E1bEjNTXmqq35+4b8lk5CqQf3VCqdK+ae2XfQNysdey1D0iGBRTIvsa8Ws+mqBPpNKovJ
QuseK0QWO11f8p8lgaNj/EpLT5Pu214G1CidEJj5eXb01XQAx4610Rtfzc/tPrdntnBubUlpMi5x
sGWF1XekryyncO/mVL2pNRonGqchcP23Lwemh53tk58+Crlo45c/p4pN7XX2rwtaVgmkUxjQfp3N
+RoZicDbb0lso/0A6XJWbK9Tehv/zLiwXt7xl7HQeY5lYziE/eebSmEzSsEGrbGq9n66AVSFe/2/
Ee6r0vK2++KNmmRVv6/IMIt1b6QxhKR9UOLhtCCB+8bmrqoE5yQpFK2zXIjHjFPvapIBoGy/qFfa
5JMf16U5vNccR7mngsvrTHbVqI6ipbnq1CF2eKLvCnicRlNBzfmWJNzSZk/9OweCKvQia4XOItiH
s41qeNT0ZjNzdJQg0qTKaZ0SwJ0ojaMs5RQvg79SvLoZ80NMWwfY30QtSVgkdMY1S/cr3Wki7s5K
8TPuOAddk47enX4Q0zsljFtw3Lw0oMX8uz2jpZQ0cU+dwpDKR8Gmpr9h7q8SP/jdc7NR/fQTt6Jy
1IrCRYEPxpm5O3UuQ0Iaw4p0BpiDafHbf3TK8C1EbRV6ShfSNSy1R204Pno9h0zuSSrC37NIKb2y
8R6OXtrdzFIH6dQlUI9VZAMri8kn0sdy6OaDs5YzZGsWKGM0vikbRjF4HNHnOTShkwdTQbz34r8c
wpuJbYCc/FOFUHaBWXview6xytqiI5LXe3qDb9LMsRO/UPhgXRRjjFgdaveVgi7UllS6Ua/2CUwO
LwiYD5fNE5H6NLI9yLFFJflbwBiMkhRht8MY88/DZbCpkx6DPvO2lMb57XAGFu8/L/LC9jfFZue5
fd8k3BsSaGGLGE1Px2VAHTXReiEjZb51pZJm+5fORBR3MhojGnEiwXv+NMaBjfzYin9xTPMu7QNu
yaMOAORv4hxNh+sFzbCsbwFliuWXwoBljvKrzkIff2X3DTtv+28bO7Z+MhxpFJyOvJM96t6iL/UQ
1lJ7MDPrPQ/1Dmtm78baTpFAbwApUlX0/Dv/LKb6A0Hnp6W6LPKJML+6P6KoAJ1LKMuV+ag97c4p
Le2+IlUTRo4w0j2qJ/PnOiksyU6/AXgm69BG0LMIHVQ127E7xjQqfNPJgZPKMkLb7E3rnwIdLJbb
Hi7t25uH2EfJZvLVkhsjZD2oyEpydXigthak4EiewV0HrFkajuUPjj/mBCJYs4YwMRZwab1DcdIl
Z/i/FkqYXtvNDrjvyW8qXqCjIDTmAmxEEgVnJGn2kEEbP/QM2Wccdfw+v7KvJQ7RjmPymtfQgNzz
A4IMkgptdvf/lVG9E/0JmUAc/wSpeVKxAJ5KJ5NNGqD1YDZHwQzSOP6R8awi0qJxe7yJ6DoSXwxK
F5Qu3wI9X88oSuMty5TzOy6R9hEEe7+ks1W4RvwefJ86bg/+xN2Yr+FURn0mpJwJEyIRXVqB453f
dYjOYrrh6Km4/bIh+yTuY6BewpL5VfJC1f2m6wIo9JJoa8b7qDxjHDs38qnmGsvqQB8KkjN+xfa0
BZG/c6v1iO0m/GYSAiqMFuzupsM5zHt1BUEjOmHaFdWBzH3OOWls/qj9mSJnitbgEmjsNUDKZzFP
lgkN4m0NMvjTNhYGKyPrqc/oVFFB9QF3nGhbhjqvB2Q/1BuRWown/hXFT5yWpFJAhgwO0TkNavIx
OfQL21PsTdKjsKiwzK4oJFucvi7DLWszUXocYHYg9gqIjGFUlbsIzfSFcfNeebh/HEGOE3GELLCK
AAnOeOWA0MWkzMkmb0RKjgsdgW8hUP1nuAgx9nbi6LXLbQdocMLY7xLAVimI8WQ+xYfHDygzsOBf
NnaSl/77k8XBj8vtGsaY94dmBwTNFYjSRbXn79R7QasHam9aO4ZjXBso12b5P9JcgmpkvckJu93n
iqJ7lLfJyFpj9j4sfWDIpMBOE1WQ5KjUbDz9SK0E4rjgLcqAwMQkYX/xRJyhkBZyQ36R6P7/HxGz
MNNj1YuN79KYf7CX+az3JzXc+1kiQX5Ec9iBSsrAt3AYc6M6CtFcvUqr2Ss5W4RS1S0h3CagbAb8
nEhZGwjY02Un6CW67ySDuBVP6aykAcbM7P7Cj4qXZbkIbYRltkV2MyCBZKpgclFDQTtndz65AIAj
doZsc6vPDQ8iPzVv3/fMQM46aX3hsUWWdpGdr+JrTkjJWYsbVAWU05Kv0qAfMxI1IkDgg3nGWfgR
tT/97i83BZl+nzH002YYnc6FJf2g+N0KxFQFUQERAPwRXtNur12CYU8YE+qfkRQXIjp9ISreJ/GT
7tiGxfVfEkHYtd7F7TECQjUKwfBeC8rbC+7mMyS9n6iL11dFUVYxQe49mZxeZQUZyUBtELJJwr8J
6d1aCVDjiQ9rBf8lk4OxRxq6lTRdYEuAZCKpbNCF5KhstuQP+/YXLrlhcZTrLXKhNV2ImMHGFW+d
eWbFbiwsUaXEl+SwqpMOwN98+ZnNV/34RsLkyQ+9tEWCQoQBSnoFO39L4/5e3VRmJIMeQ+rPLVhE
VNBqM7bY0kOxBJavuehxUtVAgvksuPupFHdikSPE+UEyf88U4IUMX7B1hQlbflNwsTD1lFNFBTpq
mdOUfdfMWDLEMjADAbnp2WfdrxAn0/Z5w9/3IHybmyWFqzXgoYSLFVV9J+5XC0/wTpAhiUw0AD6G
Fv0C+ueHLgkJa1P/fJ5A6nAjG4Cr1/bG/1JjCA8MA8+0KP9FNM9D16uq+hGSrLYmpxWJ+hfrZjPn
ljDLb/cSiRmcx8tSs7370CLTbb7KSR69Fjxc9btrdjD9La0Mo4PbzhNBB6RKkj1gDPlCN46rTJrr
eHFvbGOizfH3SxhenG3CU1PBLJCLPpWsz9XJWQP6yOkyD3m+GdLr2G6xhG1g2KVqbv1rmBY6XevF
4Auz4H49lUEFprKX76JFWjCsHsnB/c3hAIafTWOuTt1GD6gRR6bROIXzd6TKOc/3MEGz47LXdn/Z
kZv+uIgxvNgvtkcK34+vSl9X+VJ2seaofJfXUfiZv103kmRxQ5J++R4yDaPaWYdhj2mDWQMMAy/O
y4A4FhedYDGSoca5r1TlqKVscrMGRKx/Fmc802Q6iUozdvLoF0D3lzqOlsRYp9raBjqpa/me6D7V
ejOfly+J+EtNKycUZAa6UhZfBZSZn46CBFWIGCbQeYB0lPO9HZLv2VH/PljnSTXjLX3kNLvrfwny
yk+vKxnNIBKh/BbvyCR7cPy7NMad5XuZKDUc5xpuGqFjrQA+WDwGCMUdJ2A3zdY6kZkIWB1kcIPB
+gF/+k/lPxr6tZj8WVWpRT25SzxhmvuP3JdXhtJqHc9tPebMucOcXftQF3N2nOidvGv5Cdn2xXUd
8EyOwfIAqltO2dctDzszmf5v/ebquvsij13gLIiOR7f70mfLVVsV/hpk6BeIvudTTKYlOJzRSIxj
jjSh5orepNDAt8toBk6DMAg3apMa9A1HKIASmH+o1yLUoAU33X132ODUSxSYqBRJQqw2MA6jh60Q
Iyd9/0ngONpa+AuZ4+umJn/SPVln3Gl8H+ETPeud6PluFQogJq0ed1YdGmeYdbqhiqrYmP9fSlJ+
kbNpYwczbEszNzhS1vlRS/AmPHaFDpQKpTTfCZeSyMBaL0Q7/52NOIW0DCkfCrYIWklssPzZyL6k
hh4apUjk8evBmtgISm+j2hnG8OdZugoIwH1pnBBFGUOg823ihurS8kWP3R8licVMl1COIGSiKTXa
ZhA5CsIA3RHvI1jz69kVhtE/kib2Vmq8SCBC7FK2Y/wPogRbulEnj4ZVDaZJ70BLxIsFYP8u1vL/
0Tq1jdogoTXNxx+YOWMrqTVv8dQQycFWpACLCBsUsdz0ZlKHOygYJSpmuBVrS4zRsn+Z2N8MyxwG
KENDbSH0JSEzeN+nYzHuAvOYJhjprsAlIUTyaO62d0WNip2KmdbpxsfzXIThqw52ebI/Ids0KcoW
krijWbkQK/b3zXGzkng4tNgzbexNmjZj1RJ58xzllfSTuZgyQ4of/6pDZhVbH0qfxALS29XjEpQS
p0IRHPrYaX/f+pllQa4No6nHfmab/XgR5ZvcM47zg5pYr6g5wZjc0274eRem6Op4QgqynHvWke6p
YJzPESOCxjBhu9+pU1wn2IFE0mHfV2BjISOYBiwRrM61Yg68RAHofIpARywje3f07eN895AkRueW
2SiveR+azTvWHv2OM8GVFEMqU0h4tnaEga59pH6DTvNoWka+0BCjauJe8HUOHDfr/pinHL3wInju
R6mMQkRvl/IbNaaP3Nlu6bgydon/bwd3PREiDBXXBsuvXa9Nw5d54FqXTIj9MMZq7BA2JyV5Wy+2
Nx6jJAADjsxVwp+4rpF1pgQQBHn2ZlbjdoXvLt0eHjd0/vK/3YITipmQ9W0AdFJo8byr5htaKb9u
Z633U3nvyEoPGaAE7vEj7X79S/To+dgQsGLY9GHKztMz0W97u6/D7m1CnNs7enMrVfEvPGlZxSAX
r2zXx3u8cGd2Rx21Oi7AAm0/R7x1iOILCAD6yIG7JA/7HQbADR0Lsmt+v0Bv/KZs9SG3TSZw7bdi
dfMxG1ntruVcwZ8PY46ZMBMrkgjzJgmYHsIkXbX8u8hzt5iVWBfkYTH6FPFOo83JdOXywnBZmt3W
rVpogjZns/p1l+jZ1c6uoAwncQ/6pJuRXTIcYoXZe2Ix2n84GWGrFU4mVyXSfkBw7gTb+HNvD3Vh
oDU4PHTxsQxHzt7PgAJrz6zQpID8qyU7j+qA/XxI/ANfJSTrTP7fL3xHo8asb5fRs3gEKuUY7pIN
+McmvIYegcyyVj3CQCVN1XEj82wqKme10rXdnaKwF9EQF/EgZlu2MDYxWe5WntMeliYPDg9i85mE
rzU7C33RWAgeXUOGmft+0kERiVLDVveXlTEFb9Zvp5W2D8tlxXVd6r+/JHPDEk9yNkwchoUPjpPJ
oT3acsucrThnt9Qf9iiDK0/L4v9pFcoD/5EsXqRN3XQESv0f91MEWo3P2vLUlR/jazpjmJ+KnkvF
LbpureX4F/Ojw0+Spzi7FX/3Eo5y1bfxlP/DWjxylcAz8GjEmxaSdSRi8dBfRIQ9PnzehJBqIncb
oosKR3THWXniVEBw1TPSZjpLZ74N0CcOYjiQ/vnS60yrrjg8joa4BPtahi8cL15ystwq5AV4PTBG
pctHWYnexEpxWBsfkEhew7g437zDvslNxxLMfethxkcrZXk5dF7rwsPuOAdgBZymnM5XQgwsmEp+
xYK9KIpNSUqBg/CracGACyDAjrKntg+oaIPPVyfKXnq2FKH367eUHxul869ah5iBr7x0lLhj5ZSR
zT3wXUewV8BGEh7r4/oSdYa1AcVVbU6W0pExKw4AKSCu8rBBAop7pkmoU5r29mtRf3GpDb2nP9bK
3RvVkJOIymxcnUbJcekbfWLxe03ughydl/+UywQGrOMrFl5K04BGFj/5KaDZa3EFq19Q9KFCbAzx
ZvvcuX6i12Q4kgYPTmhegGb7VAM0g3vQgXHN0UkPfAk8nJItRsMEieFtzfx3RXU4NzINKEN/4Yjl
biHvGwj+vXibE+6pM2Aob/XJO+Va7cpDQIJaY8B3wlFviYduhw0uKzT1+7KnpPdGVa6NDCBep94P
yCHiVKUlF8eZvx5voJ9Lyoulq+t0xfJWhfetIKo23XqmmCAdZPr64Tkp7ts7f2sZOS1H9NwnSoHv
cQy6Xq7EsvIUOQ4FkETTitU3PVsSXAI3om881ty3ujO7X0CtsZH+/iGf3RKEcVp59G+/Zer/ceDD
XIVRRQDhGjOlMYflIAarBMEiv0eudbULb/5TJMoztUOm/a6zLOaX7Sif1We1NgMLExO7R73RqYhh
MgDZhkZ576n0JyTVnmTKm5Miq1KtlcxGLaGrPIyu8ZJf8BcmJMUoxO5H8632cDrEt3u7791hID1I
ui4WbheHeYFHYRw1TufRG0tdQq26dk7DaX90yzA5wiMkpKphzz1fu6JNxwZiDiT8/sxIFNi+Sxx+
sApdU8unUJOapAj84yLNepssY7AjXHzDAVJZnUJkl5ss8VKgh9NsHfL1hnsO4/fXrgK1N7rEzdPU
m55b15DEqVHAJmif3IOeIcuxCHhX7CDZcGLEvPLkVCtmd0Cc7897VxEV+WHoiLv5Zwa2TupNyh0f
A2TAeEUv1Od2B38kNHkYrreWxDsDGlN0cGFOM6x9VWzw1Uhy30WaQxGQu0uJ/k0w5JQb/+1Rvm+U
OvL15aQzpmHfvfuzNGFoTXMGG6ubOa+uWDrnL8rklD3+iiqIj1C0OpafLUGdT6JKjEKKDnjGBMkU
rTqiQpv7hB68IA9+SkAuoZaj5PTHEcZsVl3aifi5v+nPmwzivol9VWI3Hg5TIUS1qNnKloSMVyIx
qCSRti5XlB10y+ILdFsN0KTBNo6R5yDL/fFQC6EDRtTF4YLV7/K0AclNZETGPp55h+jyf8QQ+rSG
nO9hLWHeq1bpfD7nkdWEgNwv8IBbWR/r0akqVPVqMCMBgDlyzxCME13aQd0WHQCD5txpkeBLC+rr
gfe6X5YMr5TMvwPaDAnlxv5X/znHD5vQUF/zxgVjIe42VCoLQWM1z58CxgY+rR0R5hLn6m+RuNwK
YxP+I4SpDjDveASEasRh8hTjK88WUpVXXhaY1oZ29aVtC2wJtu3DlWOuf+AatuTOxKWN+yy8lwuQ
NnxT0cHEKSg01e2LIj1XU/Sbly7DtpHWmAoNEFriWTB/veoGGGtzGrMaOtpsRETpw1JS+/DfsUyD
1ALC4uUI3ldluZv+ax74PrZpanHkF1+P1SFrr21WMw6Kgzn/8i4XaHXki+w4LseDai9akp7ZMy5b
kBhDIIZkYgGiD4t3bsnIpEdTgZYbmY1VaBtc3gI8BALH2R+QTSNuEvv1pZouudNaxZJylfSVvzGQ
jNU/cjG/PUS+LcHfttpGW3fnvKRXfGUEm8mh1mSWFj/3zXwWktFprsAvjGV3Oz8i1MO12yl9UeI8
wAMNQI2CvmWnxpGivBsYMslSYjzJEixzsbZWPm4DwMhxW6jb3YxnFGpM+EMlaAGFzI8P1BjG2+rt
P3U06fGARLsNfETtY2NGwpXd9apbrdQrdGd4/wULSjI08adZ2o4R9KNHpAT3iFJY8nTI4opgxcaO
if275/+eRHkWFYQy3st7RgCm1sm4nb00H2O8kS4gxv0z8vOosAeqHWLyKqvR0JVP68UnNzZhrUh4
52ghuquHLHU60raxcNNb0K7I/kn4wck/lsVzzsMlr5hb10bBWXK8pTlTLr7xNW/Qj84pU2BJ2WDy
FupPpPuGhk2KbJ5LiYB67ZLu9KbVuRkM1UwPqLKAOZwGaWd6fySKCWcXEZaJyMyykcJV773gQ9qi
EzfZr2D+FXKKC9sLLnlPHiRl1jIv218v0M6+DaQdWXHFcRFU5GDs6/8ZhHDRIiI2QF+qneEZFYS2
Po2aQ/7o7zTdPdHP2hufbfJK1xSRUwBl6vv2DYM8i6+3FSA0Izu57qrKMw8ASsVwy1FX/mw76Coh
Z8R4vRFU+EY86d9Zlsd5i/BEGfBZX4QZl/0t/3l7I0wP9n/kY3Uvl98aIemeNEdbEOAJz37tEsVa
mj8gzj5pOdZZCX0Jqd5H991R8f/tR1dm3TeLK7WJW78JlnsDB9tpgpJh9y7MHhHpm6WuwLXCNMtb
OFZ8u/eIo+nI0JQIOhoXLu5bXl16ZJKiItXmVpKDe+LrbGcSIe7pwPpV5uHwzo4Ca3bF8A4VlfEk
WoYOlPiA+Y6v+b9ARMXCOzqxLq/IxMcgioweyjzh86MRnWA6yBoGLZDk5i5Pj3qKMboKHP5bt0tM
BtlpjH+DcGgDOMNrXcTbjZOq9fQaaqgCjjc4iC8Tc0D1bmg6X1TvufvPkVHNf5FAvchfFtFxI+wU
MaP4gpVxitVLrZMvvtPD/OMobJYFYNcmPK8upWBpnGQ86pm69rG/sf27qX8jQaUup5ojfEYl2QhP
L49jn0GbKTpfch+Uc5XU+PiTNG2Xk/14eLJrU5LjC5crQNJwTVrYawRYqPVNVwlO4zarDf9h8V/C
k9mf4pg7oGujKImBhwZntfEbksXhmpjRZVnVaMonVy+P2MriiSCslGOctmO6Sl+4GoioCLIiF1LU
qcaepClVbQfiPY3k1V4k5pnwuCCVWF1F2tk6aBxRXNVGDo8D+9AoEUjO4wBxb0/HRVk014143qlN
kRtLcIA6NhB2XmWgU7qXpbEqEvBbFPrCDN7dQ9YRP1YYpgiJOlt/uHb4kKaiFkyFS0M5on3SLeZi
1JrT5gQ+NvEHtaKvy8E1mjMJJ2YObThPHBlli3MWky+riHV3pWxQagp4S65DLMdDHwnzVB5VVVXH
Sr6H/Tir0a4t6p6751Got79S/qFXj30zMZeb1XgolJr5UXoAoeUSiXK+n+ur0Q/JWEV1lMO5saiH
VMIAkkc6JYf0jAMyQetI2y01ffWpbK6HC0YcNE7PLu/guWMQisHmqxZ8AqNzq3Ek95+oKLfDf1Z9
dk1IPRXiQD+YVGmUN7jkb1Ks6v7ZrDwkjwnNZi8+mTiKXw/GTPkv1l0LAwFyx7Xy2rFDB86NzQY3
hCmtOKJpKkORnS5kCwZxfHD+5bl/pFQgNvxcXtgFIZ80mAUxkEv3K/kWJLUWOJOWAf5CJBS8GoGH
LvZjKCAWd19q+2ijcc6rhcQXGRwup4feu+qyFExh7+3Yha1Z/jmEiBl9mLlLpwdN261hmMZM9nDS
vKcjMb55GmhtUQIltLlOYMvTd5pSlHsF0v3TkEQJGErmpcwVXTlpsn4P6m4VJBKEZ8wI6bND8i01
pBkbArhb/O9xPyPbFdJY/F28FgHUxXcwCTGWsEw+olS1fB3I2pbDKmiCQh2XPVgPVt1kdmxJUMbX
X2aR0ICzh3dIvADgxWwEbZpWjK8iaNEwGm9JeowZZITL4bMlxstHX2B35U5EWmH1FDELijdjE9Nv
DzLQcRkddXtOie092wtL6VmV4ujtvFJFcPSpocqYqqqzEiK7UiPbd+kGCeeEU+Iu/IPql+Dc+Y2j
bY9VRRKTx7jlfKk4q5o0VBW/EFoQivD5h6s1GZDKVqomK4qjst47/lIb21bXvEBlyagaNQRtTcIZ
AQY8KPDDAjoaykjhTzeXS0eSCWYPmUmeoyay3J6hVhFC8dT7f1iEFi6mcBRA9xjuf+crhcOjBngL
R3bwpdo17WrxQbJ0CMe4gz1EkEex5p57j64GT+vLIViRu60QtE6hpOm8MxLvofxsrZnhRDLose95
+vz+wNtlK0ffknDSB9QgssM707B2ftZx86SHFA3TYxiXKO5bTPdZphfr9zx73ZqhnBJnG/c/eMSj
S9qPnvlcKuEB2+c3Xhq8Ufi5nYNu7g08OnpGgU4vsum7NaBtA/CnR1f9H4xEI3fLtYs6/w/3a6BF
6QV8Oro0YkwnAKpRmPMtF89/ZqsHH+FIjtypyseOdvTHsgEbNiEbjqFR27QkeEHMz7m6zsyFWF5n
jdwF9wINipifrcEzjyfhp05z5gGzLeM6Msw4w3yIujHjlDrPVshOT92efX2i6rZKcfncbeI0avQL
JzJWNM3BmLH8wdPVoCPUbrgfQFMRQ9wRd5rkyOrBRxfbYceT2zS6u72224DgLcN02dttxIzFZdR7
NSvjfSBTc6P/Okn7qxuzy2ZU2Fw7dzrXxs8hsu0uRIOYOvgFElvN5Q35MHxzt8IgNSMeXnTYuMEJ
m2I+UTSIpB1+DtR53Nv49PZBRKma9YEPICzMDZ0UtGwHD1Z385EShZ5uEUiZY4YfNPc2aMVjnz8E
uZE8mBcqvzSia7/kP4luAvwsAL9jmJbtPJ476YcmhMWcJ6LsilrgP7Mft/x5bq+38ka1IHFeD8WH
XEUSOL9vKwkdcHJXZeKtd4Mvu724WZfq4bKtLofKDSWh7AmD3WodLWQFCEIOTDqvSJzDqn0Lyh/c
km5Ln94Sejn7YLhLjWHIw1SE7YcTUe18oeyutSNr0LmpDg8Rv3uUZOgnHLMpGASwvUiDQ/YbnJnE
Z10e5vPdZ9xA/6AYwH/4fzWaWRqxMraySIpffzPyekxuS7UOnTII6YR5jmVxWReG4d1F7aAABvRc
hC4hTM1taCLbLrsEUGlgGq+UtTSyU79kLizya5mzzf4RFnGB+YiRrWsC3KA0fuQstBtYqHj4ND1G
wxxYesXgtOR9cmwWZS+INiJbyM3mTB/BOLX2YPQBJV+i9Qu+V9/rEOfH/A6qoYrJKbcV4WeaaOT2
cIWxY0/xoLRXkY79Aj2Q6ibsodq+k6pELtnSqfDYGwVsaVWfMi5cCHnieZxUjsa2zQpLRyLktVJZ
cXr6xMsVtey9gL4lfGmTnTKPE4yyLBMEwJdaiQk1bijz9UUTuyLYnnxeY9PBKqQksQ48ziDtR/9G
NFshKOm1zGmAZsn/eLKiPkDUnS8qT5nbt+QPV30lT8j3zQNt3VCAH9gcZ06JEivS5aB6Wj/fs9uS
XmdgXNZYSeRuCV3FOhNBxRN6NfyOq5k6xnJF5ZY261IGckw0jweVfrENFhmSetu3huYfXC77E26F
BB1g+1pMppv9l1OkBHxUHfYg5MSfLIp3f2pbZRrFUZG6d8yZu/eOYEZMM/4akzkks3q1+5TQkqRG
IjomKIRql8ims8iD/J2k8cBu0tKqkySEof4bPbYFoVeHhXsCWE+jNiwuqjseyXBK3+brZgP/MW61
d+O2n6SF721wSpDWkBidnChqIP/rysfiD3l/bBJww1uwOMynAOunXN1DEGZtK14wmGmL1bAKS8T+
DkgHwCM61G5pSoaWwcov8DMU0ew1wk1ZzSNsDxungoZGYNDW2rbPgZH/QWGZdDAEZI38F50VUbOG
oGucquv3a56Dfeqa2It4Fe4ChBO6/IrK03wnZRSUlrRk5Q0WDPAsDDhDdiSI4v328LCvBBGCgKId
tQwsvkf5tbKg7QMMeF8ujfVi1rTYgfzmtHbTFPMF3monGo5AogTd2XQRYiW/X/KwIvnNc1sL99wq
5SnZUwu5Hk/TB4hdbadBuWNtaFj097S9kB9UwIFqzoKvTy+jdXFvb52ivxlQQW8iAINdbfkCDzFs
H3zl/EXzDPXppI3weV/TxXR/AQPuZjTUm+80ablykIMfBZCtZgalpTZUKVwDq6iWcvYKcgeJyr8x
2Y9wC993hurzKaj6Rba9uy76BaKS45SR9LUmg1/klbPKIpx9YktOjz3w/+OasggsjvYSZSFVeGgW
hzZ67hlUDcdtaSAQVfcQu/iSOaaCIZ54O3H2fCgpe5w6giWdWBkp/Hg6LMMb+fSAtp7BcBYXI5Q2
Y8Sw7yAIRRRK9wEcDhVmJZBRLT2DHBiP+jAW4/61kA4NGOX2VgaUC5DSJmKgF1lRRkxxgET4ZDcj
y5xPhgzmWQZ61NHapByl2/3ILY1Fr9NH/fA2VGDn+s+amsy+UfyV3mZ4OMDWrKTsdobNAr9w7yqE
EN6NPG1BJP5l+IqgymiEsSp2vCHrrggQAXYOv346I2swyqB8t+vSJyN9rl77hvNIFVnSbtoz0Haz
RIioyM4sp1bBcFT13jqG/iQ5dEQTcjyZgXQ9+2pfB5lXqj5etJ/91QSAPVE7EQnPecVjeNytMxnh
FmDBUPYM5wcguwHblUnGi0k+3mLMmQFQIEWzIaNchE/fafWNo2e3Ak8xZCvfM5CjL6LwAAkP3RXO
ZuprNIDrXBtGjWmVvnzXTB2jdU5lBdI0hwIkta+qCyLlAAx9yctH21Fjkr3ChSZmUfgVWEt37sjj
fxkytur5hTggF4sHKPEbL8KAqR3ATeJgaP7VxfQp7iGn29zUQbR0734yPD+9rP2kV22xgNrpDX1X
zk5MZdN6/gYjcQ11jMpsJHi2jfx4aSm8mOdPSMHXd62BslwbpslTbiNbVllDNP7/yGnF5tCgB6W4
L7lP5CimbusDG1vf3FGKThO2QHljwaJ6ZtDb9VbQtLRYo9dGvBpXPhBlHVT/IxMuElCePKY64GX9
ryA9oeJfb/uY4Y4MlTYTJPOUFxgc+mNIeTmIMFaQ/IVnv3xUVcp+A3vdFctNZ+rPR1pStjK/3m1w
nZwaG+JGsZZks3Gmnolp/KkDyx+tWWXZhKbIUEk9Mh7gEHlb3JTzk/V63pwiKQ4FUAdmKEEZKf6c
/TKAn3y6gCYjHxTj0GVP+//SzDRXgspIIbY6c1mYPe0uZVpMXmNKmLiW6/XG7wEeAxef0K0+huId
/h8ZjTTAQCpvgYecxgrPjM/iy4RtLkk9wwb+6ZUtW9l1Zs94mW7L1Yt4B4Fa+U1c3gGkojERA4O3
MelDCuY7BR/yb+6NuPRCOAcOgS9V3IeDMp0CmOGGeVNA6+8I6L7wcWrNYnKPHEUBVOpQ7mq/CGGh
3isKESIVt731mCCK60O9Yy/pf7XMnIfdVKTU9Ew4G3xS0AIaRZgw9hXztq4AY+RaQ8Mh6Q7MSnIV
ybZC9MUF6/fpTrdI6VMCRDiwhxumR5N5ewVzMkDsdqnvGFHPTPt51dA3nHFvF8GSDQLVnfIuNBQK
9gxwuCbGjj6MIwpgDo+QMCUwVhIvywYtLB0B6WmAt179qerZd47E/WCHM5RAZsETdzSf2oDVFrXZ
7MCXO4MFjZ7uYh80xpTN++U095dGYdRAJReyhDfBSa9kWzQURxGl4rKQgA6+BhbqhRTn6ZooNsAW
gzULI+nbkfhy330GfIP7LrniXKTtKcqyg2eS64DXQKX8w4WH9GjTKIgiep5UyCa1HuEi9xSIikh7
upEiZWiomJpTJM2TGyPcNTR/hU/b6IQ8Zzc3PytXJx9/UdL+/7xknSoXAvmz8rlSmPhf9jAd5biK
eqFEO5v0DgRGuNboamxerEZUOER3lZjqLG85cmcVfCzNOXJXwQDLbbkCWjn4UH7/yqb2RqdlzvmB
4/vW0f4Ed6eAZFm+xHpq4GBqpezd8n4NtVzbxtofMoFh7Beh8UqAAmX391j/G/qts+uYJkbFwazl
lGIW9+B1FIS4SdBuqwuzOTqYhF84BeJU5iCDKPmwyLM07AInK/OIpFI/MQ4CZTsrPMl5yKR85m0s
aIuoZiWz4vPoearkm6bwu1V/3ulPFDjCHT2/Dke7/KcNTHqRrCFRj45c999WeZ/jheK8ASqK4vA9
bk6qBTpiQ7qpdCevqgtxGcWdoKzF1QWoVsh3wXEbP+8tc0L0Wt11UYuj4+aOEMbtZdZeZ5t6UsCO
e1ZtZSfAL6mRB59Fc/YgfClEvPUDyuLczfKp9Dysj9Q0kjDh0eYx7fYzZZ1A7IuRZgawXcGOtk+J
RH7TSra0RuOPc8+3fYh8FIgZgp7GvSZKI7jZGIEH7SJzBPZXnrYvz0L+4rJVS60Tb3RaBL4J5y/8
OvWbda+ELnU8iongANrwEZKuRvy3Jxszoq7x56pHtyWMZwJI/gh2S9EFFIrVt4RaJbG83IvmM4bP
u7kps1vrPZq6AoCl4k5HmD9tfrX+FYCwBDHDuO8dMu/FOphQK+duC5zla9lZKdwAZc1iXrxP5jiA
apr++jDoP9PvhtgnWS+aZovRZXxKSY3KVgWhKX4qIF6Bu7KPdXOkJGRD7d2kSW9/j8gpmhcea9z4
66A1Mxbr64E2IIgJhV3weGTgt5w1zp0FQpfZh4Xse8BAYU0UB23Ys1hK8wlpFp2jcrUPrs1VwryH
GVhwtBgwJZCYlDejOIv/L2Sl0s6vur2ZKkirzbu8OjB/BSBapypptiNDv95u2DImeb3vzd+88w+z
0+6SWwlN26bKS3KHyDTxuYPHMsTFejSoNWogLoCoNQK+8Dl3shIDLwkQ8J+ZTEhBgGTf5qAVhYEi
PGLNzttlFuRD/0e+3BXj3pxjkpkZt8yjUeflGzZwbQjpTJE8YMpTs96XbQfdcj7T1nON63DppX1z
XzWcjApSk3cUaPpmJyHDqELCOuINqKq/GS4jfNPIBpV9AgQWOFuy9+EzEbH2dySgCu4miLvODbdU
4UFxe3HtsKFQxYd0P/qKEkLw5tKwr0EztJ99fCMz62YBznmCwCCxFQBBC4zFtltD5pG0al6fufeg
5byljZ/8bPCQLfPubL8WlqgwTfIe1+ccEO5DqAUGZ5x3VgZLHOoA5H3oLuDBdQ0RjFXshAQRI8Fo
IWOEpdOMoUr8hpALFr8YNddA2KhhBjvmbrwtpd+Pw6ZOcWBXIwlVqZmrQj64W7LWedWQiLCgu39t
GXWrlT69u7VjqjX+r4rEIEUDb8BYDuHQejsnFgSFB7/+3UT3iubss/IUB5a09gOnXrLyMfyb7iTi
JZJFLaPp5Mxl3Zu6vajedGo826w0zmvCdwIMZyXP3Q6+0VUOyeXxGj6G6bKcwQJvyvGrySmrfBX0
htS93jl3J48J26p0OXmvsus2cAo2pmLVCPOBpnY5SDXMwfncp9F+2M0JMqWVa49GGSuwIZy8omK7
Q7qvRq5p192BIUgX6LZOHjsQfc2GURRlehOvzvcMfX8oGcN10rO71v/gayMOMsysslD1PGC4UOje
+uaJWgNlleUewI36rem6rNsTDW4VqHCgaid+6Yw7Zq9usg7/bf9QU9JhcmDiR+QVk0nP9bd2f1HG
vSg7cqECapaUdlKN9U5qlD/Jx+RtvFy+i6lOTleaGqY0r4jheYL6SwGnMWhAPeTY5vXMoV4YeHrl
t1YxHyyuLA2j5BFAG9V3HR0tYx8uXGS3wxkwVG8diu9KbytM5UOSa/sl+moUYatokyCaBYboEh1a
r1QJHjzgeyYTJTJD+vEEl8G6Qicqbc97L7oxixPyDAb8y5R+eEPqutcmF4J3F1zyQCC/14x7U0kc
x8rj10x60pZX1PjV8xFJmjWRbnDpcR3KUSkFe8ZuCWlosQSzHiqW9f6iM10t2DmLZY4qoGd09gkR
ATDG/e5XXcNnqP6xXnAc63cUtMSjzhLOyL+ezaBn4akiQIaxv2iN+cI2s+mhz+ulM+tPkW8a5hB9
99GniclS5pY/71Of0dDP3FMudFktDvrqaFzYUOicU8kNvVxwfIvTG0aWYXuycYge+Yhp855YplK/
XNRpi4yRSJ+OMjcsb7PCdmOybak9MW7P7gkLPmKQFfSvpiTRO4AKglGTYJsBDX8zlOLHG7VHIxmK
7mQ+EjRqaoHvXCWtRE6UpwFmHJDZW6CEuszzXVaIkFbwjY9rDvC7fUAGH0eKLEcZRKKh9pkeLpNq
I8zcxsLbs2qbVbyJQZAuW4h3dY9+R5bSzf8RzmQdhQQqcS1Pb7tQK1plwnjIABmIAkIP5Zp9W9z2
QSoUBAtS8SceRFRF4XpHotTS3hQfrnsBNkCHoDXUbH0UsHmzExeRvOu/zKiRGP8cWsKy23kthQ3X
OfgfyFla4Jgt54SjNvaConwA/CXs15ngrMwO49ylFD5G+cX/ZB6JwaRBjp9htKOv3uGAhDBECpBW
TCWgsowzlRBLfoebdNheWFF42r8qXb6E/Y2oRkLbQ2UJ45PM1TluetkREhknF2aixHRbRaqU6BMr
HOYDtE9MxXQdyszlnaJODPtWf1wKm3CYwKonvSE47lHcneHT+oBQ3687WdzadgVXzU819ANc+6wz
+VwLmTwcmAm6UyjNcuqK4jWJGAwq7Kf1ycBL1mnHDdvbcAWc1anPZmSg1Qut8MNshBV+x8Zy2x6F
Nk+6lP/tXw7mmGvcKPRWqQ9nC4iu3N654P5VHLPc4M96RelbgDCTa/1BtYTQcQPtGpmtwTDfh4IP
T5z5HC1aI/aj236ETa2dmMrDlYr/oP2FEqZsLDGvX4pSa5tUeB66HqQxa5LwewsLD+9fKsCBXBZk
eCAcT+iZn9gvchGRwVCzxwnCa7C3k8jSgf+P8fPwgWmG/D99DrXHUSFfb/guze+lsk9BRq0FR9im
GRhiL4E/ZszNYMN8alLlJu2NPZO1lsu1ztewhnd3spsDrWTTYb5y25nGgX+h3M4Dl0ttEJuVGxS0
SFS8EzTk+Um6ptfIHRfEARYdTSqXfu4pAP3i3ly6LaRGXTLCSIqWqJkEaQy9jjHkUhrSVNEI2sLS
ZHfnNMvz5AaI5/vL/KVOxRxDqWxgGGP5HnSQYYt08tU7Kcy5j2xajgomJFVrC9ocoB3NoaWOe5IA
KZsNwDR6wN9f2HCkcc+tgn+0xaAFI8pCUzoDAxNbCaCJENZNp64MB33JfaAx21GmpFhQ/rwUXw8m
UnW5k0BBaJXDtZmnf7lE6oA1NTmo4Gawq6z9lBtRFl5OyzTGhsUJvWbuFNYtxywtgUL7RphbBJfC
lHM1hLduz6sIJiXoYxmaoYRjeB3jCtz4JeeG+T76RbxzVLHY1bzXpQknLuVfeA2IT0PRFebONNA8
wl6VFCgaAd0XKRZFRmFMcdEQ/U2MIWuI7vSFuj6YbJUcGfei2/T5+zTB1lkgjYaEEqUicQUqNa6P
zC5ZwxgbZ+b/xcLGpQO0WcJWKEtSKIABq9c9qp/g3+GgnWyJ0V7WalY+Oh0tx1fVjOvOyAzVbwsm
foztylEj7MLM2g5pDaC1ckRADj+zKMjSLJqycgpi5Z/CFhdePU+im4Z1USawz843mw+kUSK6BKED
FOuQBDMyHFGJxAyYrh2gue2LgJFGWZ74XEaOwIvl2LADKTjqnmoSN9RRMRM5igKx/YnJtqyNSYJr
rFgZBvvAFjUsGs9w0NdZ58NZos1EYzy69EXOhy04d/tUe1PUHQCKL+njcqH71sDE+pxtcr6/7nVv
feGYpqKQVSTyBNxSOjtCmMvGwm+ipqIvCp0Yj4l+xKwdq7i0bbEmAKvkp4N09H2chki0IqSS6BGY
5Ss9lczIIfx2C6gaU4Azcw6L2cAqFPUbG4Q+UFJgW9qmhwX4xTHb1wyC5mLfuMD8PJUgEug78bdh
lsVZA/b6gSYCY2uD8MGOgMRz5OZ3qgb9MFnkf3UnswpqYeo/VKS2jLUqzzs48j0yzhCTuR1vXTA5
E98GLJmXMYEryuuLVRJ2uCGmNAXDG6RSm3lZiWY2RTLKsR1pK8zwI+CWNdSU2b9GqlVnfviFNV5l
PT3Lcs/2unAHYsojzMzBMe9qpMVYaftJzSgZ8u2abvBWjxFu1emUrS6vcENjSiQxLtjj4ylAUBdQ
tPwpT08//6m+K0lXQLGkxXhAlyZ3e1YfLZdSpu6m3WibyyD+NQ6rDktii8qHouyb79gRtv4Kdksv
DiBRn5XxsN+GLTVB6deWcvJ2M6A7w6LZh5jM05hIKGuueh48FuCACPEZnQTGSlHw9VNaBXZjCPEH
+uURTg+0liI40kN0QmJDxJ+nbi5Ukqk5k2afZfafE0bb21r2NcyQWzQEk6LANmcxYcN6kidWiYFd
l3FaQcjOk8NO6XWDZ3pIaI0P56h2Arq5qR1hBRqYthvS6peNzcxfLyKR5kzq7kdy10TBZU3VaqbD
ugzYGC90OlnY66e4cRUpz4jQcxHbgVSYmVGa2YMoOb/c9pH5uV/CujuNoq1nYu3bhomIF/jFU5/G
nTBlxRScg8DfRg86ecvhY8faLt1mTHql8PDxAyvRnZkBzT981JforGorFccoVI1Rl2YpT71rlYRy
pQg1TBO/xMW/IonEZaz69GSiKQfFqYILtKxpiY/AzuWWcK+1UzqzsNp9I7vkpyZTigAT3SpurvXe
+wDQaqTk7V7WZ1T5VHCvQYU07Xp9OucVps/I9YEhVkWdtHvwBk9Vkj727DRo7Gcqv5lO0ENED5uX
83GBUI9N36kb85w+xifAj4PbA7x7W49wgt6SBKVilqGjaM0pGGpAyh010vXLB+Cn3j9fMDlhSCuu
gRRfsNW9EfXXOOY3q3DL298+RVFeUyxv7Llmzo5fOb42ah6nN+hS2ZZ/6y8WNivI83nFrnfjzlwm
FeZkN1CKcuvvFqjuqYSwrp5NziWh23pKEmQXqKHXmrn2aecwxWd+UAls6FYaxikZYMkprTIvGeB7
/EHcJ0Cey7mZB3ceJyDmP7wl/0j8nIegXOt2ZFNC3vSJjBxPYEwPIjqi8ZPtFaOdlkiC2aJfQBYY
cJJKVTu2hCiwDeqyrtzNV2GywHDkjfjkuw/eQhGW2kQJgmgoSBAP9lFll0VbAo+xwS0W9creIcQX
7hoX/hJUsAVZZcD5aKtrrAg25TSolWHnKrbaocJOdGbxPSk9vwUxQqXywJbKPgWeALwsm/KdOUpz
0z8t8ou+CXY7PuO5EHZhx4RhnutXfRHJqY3v0YBOaXnbDyZA0tHObbjWbAp457KJKjMCYRCQcouI
OZAyqYn/LHe1nwUMn/DOhNX77oX2NZ2f+yz2t2buGNMookbFdgrYKEJsalrcIeN3jw+Mgo0JEns6
DM5rYVviN3a7Ri82HXPeSUNk8/Z9v0AEF09zwmN3sNj9BNGv2oR4S0xy2uPycof5YdlEhuqM440O
zSYr1X7i6fmtwGG3/29T1bkXXvyHH/Uy503pOx0hGjI1w9/Qs+N3GeDcWFDfkrc0tZymiap2pexu
c6xuWiy2gwWgQlXTjiOEeLHDQ8EYKI1LohwWCThXTg/p3sfGTp+0YQtE240XF00J86cib9mwPpQ9
epFuSzqG171iM+Ge1Y8YuBlSjFhPwCdsBLcOcw5jvV12KnqsUVMKDPtfT+0t1ujEPp3s3bh21wje
aBvJxNTzUnxuIcwYWz24fKGJDYhZxIh5624dsB5D9PtbSlMk55FgQ/nP6A8vb3N0qArG21BrBrCz
P8gI6QctGcceV0E95xJ3d0OFnjke/TR0UojgVGWaWeCZUcjhyHEGHcDpXGoFGBuby8Ll+5B6g7Zu
qQJvlfwy45YwwUvKwdPfaCDQ07pfF90fM61CYgdiRn6UT5a6e5qEPYyyEtZPqLim0b/bLOToo34O
+zt9GZa4SokkU7IWc8Lt9VUVg6vABAge5NGmCyXvCgkb4u3aZ79L2EDm1gPdLRDQYS5I5v4JnTOx
k9kFJVKrxB6Rjl36ptzRgJYgrlQcn1yW71dYe5u/37hJW3N+lMpotqAWaFU4vacK6RIOQyvVDOyD
gmWv1F8+Q46hd2zdQjliInc09uPGZHKFtSWMzLIfILiSm2dWAbKkYQikCtVMaU2Frm/7NnmPa3Be
HySg1p2974hRFkci1Bz+0AZSy/2e1eEs/TbwGszsfUIsjeK2JLRLuthSe7mTOXplWu+vXBOVida8
vYhmv4T0AFLuBMzqbOVMCdlNsAyDsrqrB0qIflQUDykfQf6b5lrgd+BxYBvTzNNnwNtV31j3ZqoB
HUih4IHaU5L/AK4ryQP3tjMIodOfTYBC+Rlk5lsAiHeqwV0sQvvkXROm4W3F/qkge5PP1FPitl1h
n8TzaSTzcr/qfDexHhEj+TFjr54pZLb3vI6Cwb9sjo6/LDL/RWO5sFw7qdsAHeMxyNiCWoHk/PrL
F/kdj4fYp9k9oh9uAN34rdBsGsPk1UtqQOiOa7Yx8QWAUKTUGv8joFf9tYO2CZ6VLRf8iyphtb6K
wRhy60ELwZcdeTtFakA2ivXa99ylcloXku89aK1HeFt5r7g42d59xfOrJJqzeEavuOVuHTQXJvbs
Yd2GDuqTZMO0WVvyvXevC8Jymmh02EGn8C3I5iYD9Hu0fEd9tLXduuA0GojwgFF/FxuW8YRoSqAv
BiJBLnkixaUD9rx+ehEnUvIpJREvdCc6JuN0XgO/rGLjEc7kdQJmVsXneXPeXKV3vSPWYvQeFDp5
bZPVqUFp/jwxucuT77KqS1eYHCm2gSGleoJMVwa+BJUlTjgcvsL5nFAbagkQ91ygGyYShn42/A1S
zd9PruCenBY66oamGaeEqOzbA2pb7HNpgdAPRHvh8XWETAfGUxiNlbFJIklyTHYhY8W5G8y0FlzA
i3d2YJNtqpYjpIlUdX/ktummeIJNxhPgzrpfakz/z+Gl/OZcAqp81bD/OJyvazWnUnd8684cs1oE
aOuoPNonrk6rKt4IZj/86Oo1F0pKRIpZ4XPQxvh13diCf999rADdKDd7TpgKXcJDKKHnSRjzx8R0
Xf0dLrpNuYma1Lfr9kB1rQTZ0rUcnY21MCEjUpSrzv8rLha0EalvcXeu9spszetX7cge3IuuS0B6
llNg6HNnoHvMb7W3NV8OMP5ADqedgZiNJSKIGVsc2EpAO8F/XrPgpGqaVm7E6G1GTyAk6qRc25Fg
px3lx4tCUdluW5LWqyTK5FmKCqQR4eUka2e7HC5mHbXdKH5SmtT0q8+zbex250+dcDowmBnWcZVy
jaUXG93ikr9Yy9iY6/iR6/ZG0neZgjc8Cw19WWRecrPKN55KC1Z2v2FfwTUlc2hxofJ2ZyoDiZZ+
OxXCbJnaAsaULeASjjLFxzUK+LHRRuiLWYgvO/v1ukghsZkTW78eC4PvT+VfLRZsBspC9Sz0aALN
eQXEYYxvPF8LugpRGjDuQ1zMHh/e6/n0RFNEHO1oakGa6cUzWXXndq6SBQdLWbrBK22IkagoqYTB
0uZcQR3pS9LN/imEO96zg7SbDjkkJv79tCmnpzKkM86/9eNQnUvLNxkVlH/OnmdObbcUr1brvfrz
qUCIhOPJTZg/SDm5d4zNOzNf1iy+AETFSl4oH7qB40vSTZ83xM+c8QJhVTO31vI5eiVhkIbG6ntP
OYmKHqyIWUSvrUboC8XX9CDzQcLX9aj9KQ1Y2ySNof11zWsD9dpGNCyfg6yXHaziyuPvQxl6w653
XnuGCVKAGiO44JiiVjlEW3r8LfTH++Fr0hJbi8IvsJ9ktCdTpwJ39Yb4l6LsyYykFQm4In8Rik8N
hFaN4boAmz5xt/n6+EaIeWehZ9KtEQyuzNpqGFcbMvWF5tAPOojVGgry9F6NzCfKnkzOv/f9tC1z
ILzzKntTvgxYpo0MVUqFde9U8YPL33DuHHpHZXZwfx1qWysDjaLMFUGu3i0V0Rvh3OtaPVa/vFT5
JzrH7C1X6hnhs0TJ+CBX+j5/7ob9vXBHJM7CzcwCVoPRayf27xh0qc4w1PBHTH8YwKv9xluZhj5d
DjSOhknB5pcWOceQQyzEeH9EnWP1EZQ2i1Y8QU2meKUXndIDVUtX19ZgF2iCzT6FF/RYes+RZB29
LTZJQuqmbYA8qIaA/OxjBu7Oxchy4Us9ewP00/qD3/3DFCaLx8B8IoAOHxPKT1zZGHtLMjG6o0za
ilfXb3gP5h2XD+BkcD5tq+Bkq2dtECiId7VKTGu2VB2z24dtrZl2FzoHfWgAO7wC3NrqsQdKNDox
rUm81kR37p4BjOghMxEAqPIFs6zmcIPnsnQlr+SnAndAlYmAFpeRXvfbwvCH615Fx9LKH4Q2gKIo
hhDbymmFnoXlPBaV8mJqmbnTnQwtWk3aKYBKgNAXUOb1BSsBveUOoIvjkNAuqZZFvvReZp95Mwya
xEk9ERGxk0JVmQQ7tuhg9ir1CHZ+u5zTBn/WPHt977Ab9/Ltb6ZbR6jj5mCxESqXRz3oEw5uFrhn
jIEiA1qna2YK68SuZmlJTouTbq3RGK1sn0v2vAHkxBXZxgTXNkaUpM2Cu0ATpFiMrGYsd/ZtYkPb
R/FSUTWskZ21Zh452aYqjTSIG7Nz6TDFrN5LV+XOBHVXgz6SykBDUlcoSPY0XssG4GMoIfsOXtsX
bosQkhRoI1V5zDv5giXljLnMbZIAo2+dnxmFHfHIURGSYB/8ZULnFJTwY1TNnF5EPx/++x11UKfH
/bIQveb2f3h3PJco9XHNKSx3yZ9U5EvE3nq/bRwK7VGRn3dwxOmMq4t1LH2Uj2tX4F1bmwHfByW8
wgg+/c0uo5mpROJ/WstkxC3nSbnRxWUQrJwGPM0Fzi32siTy/AISw1TsLpglZz3SzyzXtGKFD7ct
Mjj4xws48s25n95Jsavyk17foRyVaw9uOkFwyT82jqI8nzXMGZa+T5Tnjs23u7dmKr7hsZ74NGLd
slzcDRo3IjcVT4nUtyUNOR+BOnxHGflPy33NTkab3CpLStb3DNMi1UnIsHM5Bn6zrbKuQv4BHs04
QQk+bA5G3H0xWuWGsVnpeYUrjL2HxeJwbVaHQjPAxPtgsSC0l2txIF3VL42MmPGtwB1oNksi5Qd2
4BuKEiarg19c7kcpM1ywKA6qauMxSI4yEvknqEpQu4qvPOf4EBRrcKMwNLSto0buogc4xwOKtaMu
DSszQX8rmJ2rlnJTQjCl0rXXpmAsDTnRzNHI5JHvS1a9aa2qHvKFrCKXjTGMIJ4EZSg+gL55jouf
NBvUwvgjhLqd+W9IBBgddL3uDlTY6W3vs4k1ZqDVNDAh+JU8JpE3PpLBaIer3Jo7HTpyX5t7UELl
o/J0Sx4/lM5jjdzrUrW8wSjj80vvXc/heYoDE9orDRe9Sjm1CDob+Rtw3nljV/Q1jGzRUfs2o44A
SshTec9IEOaIy4ArPi3+5SLqSvLZ2iYhMCdBGKz1HTyKKTR1fF9DBJKvOnCLMM8T9N7pnqGdx1n7
zg5CsV71ZYkBT5G6PIVWo4eflXBB2beNUCPGUs0yMaBb4afWjVT2zp5HehijoydD9/rRhbUy8Oua
fsJgA6hknRI1CwfXhnuP3fOovUAzc/Hn4NNswa06LoiM2JzFXwMjjtR5NUnw+GEP3yozEJedm9sM
xUQyzZrZQUpDHQU5UZGHnOFMe7duMuZD5b7pB7K6WjXpvRT8w2KlkG8Pk7qMueRQrMdfDwvvHQfG
4e3r2zvk0f3jktn+CzgY2CJxnuKPmj3fGvXOtUnHTrplKUiOral4G6QNcI8tMqkyCt15IdXeSzod
9A+uXkzdSoj2v6TIIf5Ni6mE2jY1ulVO82ODC1tSv50t1Q+9oI0JiRVXDG1XyOm0KbMhSNMFd0aK
9Y2kjSSYI5NGfuYuNkC97+U7aPBvp3UEI4lq24BxzIrLKbtWFn6zk2jHfMzCaSsZu7HX5m8wiaSI
BVu0bbzeRdsDHpFaKF80LFqqWu6ua777dPV3JCrhHEl6NaQb7FWpq3KbsV0YG3PZ9iNLrgNWh1VD
oV5zfm/VcorDEzNc5vMjt//fUoz2BscR8L+hPutRehTFijPozdD3sFFqjL9QDR/kLQ8FoEvr7uKH
Ga7Ly5QFfc1BxOoUMTJpEb2KBLTFoWa/09rLuvhbbyoUFlEWzXEfmeMWLUcrUAF4N166X4S73n9h
T2VwwwVWl+YoszBIyoCEAZmScXsmQx2KLal3OqiTglrOzEwPd+VStyWn6dFRruB2fATFyiE6wygP
DdHi5ibizpxqfYSd9Sa/f9/7tEb0DFJ/C1jqwF5SZCQgwxChr6Dn4lP4UxX4xGi/JxfdIT7TCUfw
Z3lQnFuwg2Kc9itCxr7BhzwfWTlRuY71l+pXyeRec9TK/jIXOzHor8v7t+s0xYXICQqAkHuV2riv
5Wvhu1E+yVfYBJ4x6NkZ8EOQdDoaVZAqnLa+sLawX7vW6G3FWzxhXcuvkLsrA9t9w1/ymbo3Zdko
+l45em8IftBQGhts4EdsV9JlES+V3cNw5ViI7z+OuSFkIXOA0bHaFb+O6bmS/BYEe/17O4OHTH0f
pStUvQSDO/94vEX5+Dz5mqrpu5KWdJqWD96/AcTO6c5aPFQZiRHgKK4PKoiMhZhc4CGubXlsacLa
pf2HspTS4zsh2AMh16SEENcOENS+8IRGrFG61ikY6VKNkhc6z0E86IpHYEpPvVzx9rLtIXjUgkGv
djpVTqe5Qu9s0+Xb2Gyf/288VG6vPPMoTyO0Eej1H7sQ4uhdaat/XcgkHisJm/OMXEOiVgR6OVKz
sI5GnWcfr0uFqBABuHxuKVFJpUDWYiHR7on301nvTBQnY6BZeq3HZ90t04u4B9jy6WnLFahkLUYS
+CTAml36Ug6/iNBS36lcuJW1aIMfC/Sm+mSnKd/5KpJvht8oEOPg+2A/BO0nFdroIebl9yOZpy9U
xzVhkdyYjkQQ4PEO5eLkrkdietCgZgbqVMiycy6QQ8tnYMwJrt+g4T8ycp0Rni4OMkuNBgfYUs+G
zbhiexbMlQ1EfmRboaRDftgdg+jH4oLro8B8v44U7kcQ+N9Vtd60VZdmaZQidcYzZypu++TTHEt4
KnNnDZ2Vu8HPyPp6EStbfCMk0nJ33EcjOIceqa9u4JQjXhZbTvD1k+Es2UKliBPqVFvfuuLSF2EV
PkSH8Ty7YYvy07usZx5JHe/NRJsCDcueorc+yjWNAU/fWNQNnDGlUsCyZJspUOAeNuXl4s5XU4cX
aB7fcqf1cZqXfFkt9jSIXJnJKtOuQXaVT9kTwvn+3YKfBxA/YfiRUkOXPMtqrGrnhHPo81QD1Cq+
a3r8iqfUcfhTdTj2KVapOKgje5yMsBX0WQgqhD663af0XmEnRSFuUlneWld7SCL9NMtkMQvsEbBu
pjOnpFJ52bOz5xJxzBmiwqsv1QKTAQ5HgGYuOoVDPOTjvsjXoeiNNLxoPYWCRvcuJe9rTvuthON/
G+bGgrfuMnXA/dehp/xWoqML2E9Y3GNVF0SlyRug9HUOAM+N922zktGao6fbGwDpunkpKEBayAY6
xB3uk88HtWUkKAQPn2IG5pJmV86f+ZxHRXzvA8Q5LWG6LPdWYkD5n98uBwqpY/L0msn/7hNX5XXk
B3Do0+FMax+Or6p42px9KInV1ghG7resSrGXlm3rMkuITcADk1rZQTgbyiWhHMh0oUAiRgyFt25Y
RKoJ0KjJmoE/NdwLgAlkVyW1RAtd1kw5+hCfP7djg7K/eTwRMhSNyYbW4GKBrs/cgloyUya/ttLi
MT8Uey/Z/OF6pq3+WF/5p9qhhVwJc+WLHW4xQLJ14M3hPhctBC9m3rGih6wIZ/H27sE1rdgWp4FO
MrOLJ5vG8a1iz4XwiGRssidvUkrh4oP5PDDsPUGlNO5CmYNEYBPlz1arl4OnqR08p9F19gY6wR2T
kYv+yxSbDKYfxITHEU+g2MtAqryz1sF5QT69DJMeOK7rzpkssvxsrphU+rP96M55KgiRxBo6dzJ1
MpvH6QjykqvOhNhyo8OiTe6qhBdEOLoFdehPQHWGA8CIxuIDhAEVDYFuVKrqJ3ebRHmUv7/0zy2d
qgVcZBucKil4M94fo2At9EJowdF+jUP+raZrWJFf/yJmg793om9BDGkgywLGR+2NBbQ5q26D0T0n
enX5PhI2Xpb2vU1OtQqjKpy+dBzP+XWd83WKextCSOxzpVXt4E6qfUacpFbqDsCMnt9JFhkGRODl
8SJrZifD/BRygrbhi6mS/NFMC4YhZ8RgKLWAURvqCD+23Wur4FlCMCrdAaok23hXlAl9D0HDwpnB
hLNdQDYd71iPGgZDXGasffF1wBUhWHEraFSoSfGDMW3pGfGJ18I+WKHxvxnaKm5p8aHKyH8rULmn
Yty9u0JPLX7pftrmhCn7EuVZCTpH7qnqgtrj4P1OAFUHWQjwu45rxE4SCtBDwKQhI3lkTMQntwq8
YEx/sPjnc9qvlla822Bam2bfeQzmA7BomcjXV0E4TydNfAcpaCAm0HqFLiu3MMTQa4Q1RBsfCXFg
DRRNjdhF06ibW8sdLoXahMLzH2b/Y4ON2W8eH2U8rF6KVUAd84ixdfO3YP42Cm6zsZ0OuKIhlzQ9
BByqb1T7W/FIVhXOZ2Apy4ZpqXMcW3YaKtxfVpSn6zHhRuY6GetcYhZbHP4jEK/uAEoQaWy/blJ2
7/NCBu3JevN1rJGWSeu88aEmJ7b2B0NCCcjnsPp6u3795ZMCr31nxiuhk/N0eN7DHkaTF0vt/SbF
7GRcrjIr8PwDl02p4Onf3hy++xlJRRjgWNsffkwac+fiLMUrxyOfri3xSnr1LmAyv3660Ssoob7l
R7f9EXWWaFiM+58dHx3JdQXYGLIJDXGQ0P4Jqim48PwK4TY39AESmguvKtN4PVQHln6iM0DChIC6
zi/DbF2Z/j7l8TdVdyWOvJ19kFkvD/TjTnS2xCR4j8zU2s7oNObsYQc101JGT7YjlRA/QAMx5vjL
Ju4+5zuwB397sSQYgampVm5FQTcfTMxmEQCgkTjEEt9XvzZtQpg2jo7CuoJTZU72etBoT2PNwmNd
ROjWV6ilYT/szY9Zty0q51EAT8MBrdoDECxCms0zfANooc7i1mwV/BvvEKgAL+E53qzknvroL1Mv
uq4TckOEmthYO+yctD8QK28l2wOe3dCRnj/lEQD2XDIZPYN1PnGcmC4pvrRwYFAMBB/CDdnUbcpz
1Pi+N7XWqRZowiuw6bWWMt7hu8Vxhgy4Lv4zJNH2UOVk6OMdc2w84/UGkUmEmjHafqdWZ9/IqvSZ
7NpUVL7ccJqslQyvzGHIxqAcxv1hP11XQpjKBdzdd5SoQ1EUtdxigb93owslM1ec0OMU4vFwYhC0
8gIWZyQeUNSrjoY9LgPgET3e83ppMuPfGIBp7se2cRTiS8rkNhyIvkEzpni2AZ+E5o/ppGcHMIDy
4Lwz3xoV+MRdC9nAunr9YOx5KBGgrGQ/rwY6XQx7Iw2Etj/e1sXlYhTsGhg7bziczsGF1vKQKK2u
4Z4Lh5/mGjSlKryLomsSfIWbnc8jJTtCUMUlWdsOD6iXVk+IxOaGQr/zzGw70Mv8hhDH0QZWT1u9
WgDaqCAKOApt81o/ktxqB9iuERiNZ4Ufaal2HCOEMcfRKiPTwqtBheIU/XhmsFFSJc3nAG4xtsQ3
Kh9e7cZofLEu27769j4yMFqMPjWZLcaPFgsD8IzSnMF4ID8vW5TEEbPbFpuiFRc5VwQMNTpc6/re
t2mD8c2QN2xbvKU3/4dDnfoFOcBu1Fey/ML6wJQ9ID/ujaXWGX0qZ9oYJl3RuPdf0/REI5Qe5lRx
llmvhWvgJlwv26TfCljvuIHiz+T/vvVumLMtQDZdsMzb0NDVPPBiYhed++NBwmwVxQ43PqjbGY01
1+2JvyAAFeSfshjNjo/JOgffHz4OS1DK9+lKlrtLD4fD8/HoG6S2kwuDs0z4HJt2U7nGqDsW859A
1V56SG+JlyNPtnLHcuIY6GsClh5EvN3JHJBDVyHYzp2U7apuDyhCbIqQ6R1zWOhAd6TfGQce9otb
3mcfIwbpP3M76AIrxMaU05kMPEew6uy3mmONCanOwNMS1fMOzycywV4QzSWosdZlx05j9UzEwU1L
RrWibzVIJ+2tNUkRLpPuXJGT9Qu6r+9KxBwnAUGgorrAVL8xKqGQgHfJ3neao6Fg0FxxT/dZXc49
IKGSsVDk0HV3lz72dBtncOufn3WBD5hbX2KUnjkNJn4eJMIlr5WBjxDGp//J8MmbesToqH20Q9g8
Al6nVoXamZFiYXpPYQlv50h1HyCmPcvQiFmZHYR07igJ6554A3XuBzj9Dsgl/dPdBPMVWpaVcXiJ
gOzbxwLPkrNGSzMhxIp0M8R08ZjDxqSCxkitI4KkYAoS5gL3Rt6kOEhOCzMP9qS2fj1Ajh2lR+6f
ceOP8ONfS9JdGCKfh2CNK87+paznhcs1V/qoPjOq8MWp+kqyO4ZSXgoxQ/2vJCg9seweeI+QZPKj
L0eHxL7ctZEUX+rIpm9FbtYySMk5+KtCBg0ecOmQ0noNJ2ecEm57qMqmKNWAS9my2AIo0UQ4TAH4
zETkqgtLjUk6HJexhp1GW26VjW4kD66PQQDqa0OJ1OmUVsujGHDF/urcj1e8qhQQ6fbgx7mzgHIO
XQqd5x9qwvP23f70w0IRBx1gqbaBd/LY8Yt8ibz7qZ9wBOcuEcm7XVSr7p4VeFumFLRgrGHtFT/p
4VWpmCyBby1repLT0mJILQf+c44I2agTuyZ4WpiDH8VNYFolvKFoAXT1Kzzf6uQLo17YWFaz3yjm
uZ2MV4vPvmw419Xb3EsqQxPrHEtk9Or2aY1FDKbec8tmG6Bw85JTo6/Sg07xB4Rw2F/tr0RLnKJH
OmgRkhcAn4lLvyGzAyDvH1FD5g0QWCjWnJ7EruThqKwCSRqLXkwLTfw6hdphlHMz8kRk4yuLaKk5
DHs6Qx3mDw5T880O/6R/rPgaBaW5pXYkJ6EcG26R2O04UIQHkPxLD8UCoGcIQMjJb7MO99Y2/DUJ
wyIaJJwFRO09GrGYK+eBMEh1PibD5hMIqybm+MLguhIhhW8gDXj4OHFKvhOtio0lsT8V8E5sFOyj
l6+oTbuPvPWEwKz0Vd5vHdP7fNKJtwNzHyBXw38dWh4hFlPS7AQDGxwNq+v60B1O1dDzNmBUoS9u
WZ8K4Z+zGoqHtqWIJL/OZ8I2RtWx06jOLB1x4edqHhLPdevk7JJItmfDE2IAnMmrUdxTd5w1+Zk1
KFXuYc7377NJnEZSuJnUv7+2VMNuCbCbDH/AY919ep7Zal00gnVstHPrQ+oC/XzJyk+3KzRHGkmB
0L+vpQ07wbcjDaYZC8qtSYNedS2KTYdIoxmqkBaKaCJIGJ0n7KkNUW3Y59vPozYf6Y/OHqQTK6fP
rJJXSPmyaW1qgvoZ8eeALgX1EsD0MzY7B6Rx+Cv7x1Fy1ndZCeeAouYD25/vx3VRH8y2cVN9ZwEy
dHpBfFy/6QVOePT8qepuTijcsmmVcVSszcPsOveST0dt3eh/PDSnlaMWrSkJTLrurUQKR4NZdpGG
2VP8TPH9k1Ml8AbPgh9DZJbNZWDKnmdKSNQ45xsV7+2TQNKhQg6K0ISgnJOMePQ40cKGzKU+32oy
sLyqjKqhg9G3200uoY9j7plzxQD6ANZBTrrFG5XgGYgWv30x7Uh9h5s33MIGvLMUTd4+ytd4Imt5
doR5f63ViskmBDjyuuX629PgmtIE8tz10M6Q+mnB9X+TFOCrKyboUtAuwbmUhYL5OgfBpvYy/fKY
mc3O9HQoZsn4XGIdmDaSCxwZMLAh5TI97CA48DgkGmgrcYhYtLGdVfbn+XaamT9RRCUxOdJ3IfS+
+w0QepKvGbtNBksgoPSJbSyTUFMIhvNUEMcJXEzjEj/JHt5eYGu4MqKN1YAUkASwEQYSQKOsLW54
cMgnCgh59wAdWDGPQby++ksdwmGcEiIcWSoQCw36SAk4s7+Y3CUj7X7KZs8TkRIvG2XEWTipe3Jr
VlcHSEgqyHH98Fl/dLRF7EWFiKqzZrDt/54UqrHQ0ME+z7qAF5U4ePpst9vAYkh6t40joJoaxXNs
P9WwutnqeOgJd/016EAmaIlcT4fJS6FZ/qppR1T7v/5mUcEJwCeAKI6PrgpNQbpnFA5aSxoc837w
VUe1OgVYT76vUBQ7PPrVKdgXwfbK1wYlXQ/17OwblBsQwgcD9n5uifjGelq2PeeWht4FZN7/zNPp
KVlaZYGsIEhBRorf/DRfyZG0hyqWwY2r/XHL+cBDEkUNcRCZ4Rz3sw5UlhqVcV8Xe374YfLEmYKh
1XZp+7a6xUwbXneegBXWTofloxi2JN82w3RjM+dEVuxt7ucJBxrQIblMkAA3612iqsost736jvzF
WzkQHubD1u392hztjXLUjemAM5sGdpjWpQudw99BSHvGZJnmI/pvxIkQnMvkyd1A9yFA001fxF7v
R8JQyEzExZJzFlD5S40UCgzX8qmUh87gZ4FXEb+Zhx0PT0qJY/99cxX9Tnl3veW38rKyWD4jif6U
9+oet0DGv1+Rp27iaj4T6pUSEESqRP6cVFlOrshvWpOEqLyl1FxNCvjKoS9gqkeAGyannNTuKY82
5w911bVbz3VvHYhxalTpAhg6b9Yacc+Cmf2/ZIr7/P6is2t1bQd+VAU0GSjEdDhSlWFyIAZGV65j
yxe9L/Myf4E0Aor3+PdgQQmUdFRtDwV5Wjta6eIP4xLIyABTVNSCbPyR6UHG9HTCf+jeBcpghuKq
AqpcnPZhfmWbv3aSI8rxHiUFpJSf6UZQfjxwEKvN4haxJq4kj7dw8CO4owDpwxPiCRdI3itgmK0Z
aJogn+eBqS9zRdOG3zq3cechMtaMHxFODbyak7a0GjmirdsCvLHGKzyADz+44Oy8z44y0fBY3JKm
oUR0V31E2T28V2YqWT/ju8GewTzFRYJawNx+nivrXbJZBfzAYzaxIFBOVVfdjbWT+AfRQdkAIb/N
ssJw5PJwNEDK7QyuGHqNbj5QYAUtseCrf6WD770h67K14vZs481OXrEK3C8y57NoyRnYe3kTC2Zf
9J8Dl7Nh9vBtqm2Zk6T4wTOB4mbDj5MCkEJkX3Tzr1KTkNCiXdyOxy32qTFcvwt0e+PiwexzCtOk
NuMrFNLw2yzXXIs58s8JkSs4Wd7qX9jeh0oTJZaWs5Z9eMn+0yS8Brbm1S39BBNQYJu3PmkgYBKg
tGoq/rvdTEVp8+slF1LIWmLjdaXuANcedcERkULcUIXOy73wX6UGzCVHfGtxGPq1ElnVXkg/QWVM
dXalIbtX+qTcha6bRsshLcIluy82O69MuqoZ+Tp9KvL1L9NdKMYljbKH8WwZnbtvGi91y19egMzG
TaRKN+X5Dd17zySi4tczWyPf0xQMenUtaX0nY0FemUno7iGbfolXuHohEGrWgG4FZaV4SDjqoX8P
XSNQDRXK+srmnrGTGqk7AJCN2kOk3Y66exLpkcu0SE+qv/o8wHim7KwzC/i78G5MzL1C0Ud6Xu6t
FYF43q07oi6knpRXFzoAw8YwU55dp6i1zeZSaz27qJpw0RDV0Ft7JtTWpZiBZOXu9DRfVdQC2XqL
zu4BQmIxprW5uKLKqz1j77FbY5BLEgmCgMHR2cWndBdw3iMSJejxvD0JaPCTQAXOJCGx07+y0Prj
gyF6HXDkvfCKBoF3mBsuKa40HilDv003yXqBwRe7Tof54J9klsWxFtfRiryGjkDUW3Y24PmqWDde
GS14xRanBRamgD0zHk0r3MsnGnJLaOsPkAAgLm6Zgpntu3KTG3Cjo8o0OduHVVl85vlitaqJLDfb
ei2eIW7qfTHbacxgwKasxqKntaPC4nQ0koNnvdzg5tUf3CW56faqL0PQlJDsv0TmZJWTqnogTbxV
je/tIvP4Q9vdfZqtobXXcbnNVCdH9G/nPY2cNt+2w40S1E7VfddC+F4lj5/1qxthlGbW+H3e90lr
YmoQMP032XC/Q/3VX5MoDS/dvB9+qf1OjCipH0z174XaifGb9F18ef8k4CBuwtU9Qsvo1Hy9kp4Z
7cxEGYRUrW504N9EHaIWqiRen8jS4qVXMAfvDhRTWFhAq33kDTedHmAOTeZdRnMjM3HNhsSUQYfj
e2dbwIHN5bxv12F7GpuH4JRafl/wb2ExVotfn6aBKM3GWxfuqMF0yTKeYF0salPYW9w1X+wSTX53
NURWjK87TkRNbljtCBsIohx6/8/lXZJLlSXAFLK8SksTtDU4BefVyPieSfOIeRsv0qRXgg6lZx60
igv+KA1HkWIgdwGcyuhL0te4OwC9B8XPq/+z4u992wMcXH/KqJuSIf/k59TzDVcus3Xi8TFCPAw7
8F26zAuc2n1LMhku0hGChoy0jorsdhGuN4rr+LK6mu9aC6Dp6W3sbzV+Ta/sGG+r9dTMdJokrBVQ
ZB77G5u+clI80i6vFdWMWX14vIIEU4bxssJw6EvbUIQl39THZEdbDR4+7sEluAxUiy0v7QCCNlwZ
UUHSLq4tUxqeEU9K5a1ILfcQg6HgqHP+7Kyhuix3nsspVnr1AEk1fujUcQrH1nn/a+WpAmadRQGM
fEJev7rVkNIFnR8HqAWLnTNK70fhm/G3e6sHJDUBJb2bxAnQflpK5VjCUSsJ4FQxX1AULNAmn9ND
DDVhIOfrwzSmBsiHElWgegZPqPzRawRMd/6B4Cr5foGC5sm+ztCAx5M9gTbYa/K7vWmdgKlYGaYp
u1A/V08xqhq8De0mR9IAO6PCoQMGXi9ee7mXSONU0rgS9FONsznDxFQfN1ZIf2zYPIc3JdoqCJyS
ighztajywociN7TP36vmCMcdaz+B8GwFVUltPuxyeX5zpyqPJdTmCyof3LKfybQn0wov93Btdg0y
IWHfBRFPcmPSLUZzTk8O8Unfa1i1yU2ZEOMOvjlou5N0i2wSBeB29aj82bJWuUh/QQHwdNy8qBpX
LwlhYswgd6TSBJB4JJRSwdcb/tAdqLdq13aZK4TOZMqb2O/uO1yJk0q/0dhQ4q6g4RQsyScLnO6P
lxNYWgEhC13opIOQSPd9Ro3O1wuXDrzht3p0XjvTp/L05rVC3uLQEetSBrOGG89gukzP1qmxyJpK
qX1ufjcQP7iNg2zNApHMJcaE1i8dwSga8TXSnuJEzctX2RQr9q5Q2O7UnNj6YBQBj/Flzwl8IcSI
z3Vh2elIXoM44ocO81mGxJQn8JC6taJM2GOWszg4La206OxBeGpc65rqq6GEHPUWMIHLp/FFNVIt
sUcGgD35Evvrdh/zSwMc4bXCjDOCI0yiB8Vp/7cguGytc+5+YRpWPvd4ul0qzCoLIYa5nWwFNQXx
N6VzyViYf5jikupcd64CQTV/knB2O2p4TzDXS47blD8vx5jQDlDcPfEAvcCr9qDrUW+pxAn1GtaD
/u+cfQzvD4NISrWJW0tCT6+XlrwU1z+jjrN13hO+ctaMir6yv9ceODjHD5ERgM2JlgaOAgh9KMW1
OAa3dhJ/jidR79ZkTB4mOn7FJJfKSefAFg5ASmqmPN8XikMuIpsQuvBIJKCD0V9SWbtnspEp29u8
1OnXV0DUpD51EzDtaCdBeZt4Yk9dfx2MMZHZdnXE++enHHY9bzbCA1BQoBsyEF4gKPqbUpGBN3BJ
amdZmziKAPnvvOtJN4UCLFpaOPh/H4/LZOR9csU9EmhAGPoN9n61gGwuPZMt23F19uaq3SDAzsUn
ZubQFflL3hPTSdO3HUcb2Xao9sluhoO+Y/sGGPPNgpHHSOZr0Y8wfzHEipa943WbfoE9ucjmxfY9
mMKErDjGK50cCFVwKtKSaJGRwKZrFYh2oZOVlqorOKhA0nXqlAu69LBY5auPLr6OThjkhzuB06mR
r9SolWWJhXsoPcq6BdZpZZusMdPk++rltzx9xOwp3DgBiDTnz8SIxBu0zOVHByAfXS+C6PQ8iOL3
jV0GUuwpy/V8q96FNboO4GGDtZ9ClLw+GDafXlxQ0zbsBolYpveI50Q+LSmttSZcgu4Ey63H8GaO
qc99c1DoGnR6dslLEhYE1ehkizAN25IYT9UnWvhOBJzI24ZrGH2m+sXSvRpHB/PintezJoBQ7tbe
74681GG/KFG7EsYoV/diGghR5azyTTieVjN2w72F7cQblkD/4ypv7vaZzzfFGdPNeKUndIFTERP6
GkmFv6Jl0KOhSTg4ohVXFjahOxvQy/S471Ge0C1czl60QhheBHPdQ9Lpy3slgrc6QsRlsYNB9VBc
IGdB4jpfqDqOuVkZbxBSSYH3Ah+pO+y/a5ghp3FYkp+5epD/cEzGJRwLqIl6HAHrEDhJVdgN0Lk9
jeZilKAfxTkaaMx7knrHzAR89J3n3CJbcmK12R8X8eFoT8KEvIyWD3aUwdFwSkueKjdQ1OLxxe0L
9IalkfCEd5HiMlWvNJpxUgYyvfGYdR2waD3ngvdWCHEkIdn/8A1eWxTg+D5NeCSZz84fI/yZf/Kz
OHYinaQ71NcLnViujDjudJsz4twWASEjlTSxYShDl3SveY0tN0nIV49Xskv2nZO5R/N4cCJEjTbU
gOptCBE36csJly4Sp7p2ODu0plCdXjBJiThaUbpNizNhfOI85q3GRKwyspo5r9zqtvyRGPnAdgLU
Tbvck84kMVxwGRqRlt0SW0wpHffnl085uSAv43YuaYDIb7an3EAsPHIfoo8lM94mcKub4Y+NjQ9O
01Mx/77k8TNZXSPo7sfxaYIbzy+wP3Og7HeNhxZHB5/TmbD7YTqtw6cCY0NJ672kiv/m7HcJrkOL
CN8PzwvxA22AszA2Bdilvoumx0QygOstyxtmbWCAjireCLOxWv/0FECiZUJbifIHBqNsB9WKKX/q
nw6XxsymjiY0gmsRiaFsJX/3T8TFnehLQ4nLPiTduPlIpMni1Plq2+HP2jFetFH+BIqEVnjQmYiq
Fx2GgMlajql89/ArsM25lRhPVSJZlcLccWXZsFtJ0XMaHmGvZ7rpS9q1Q0+tB2JXat5PBxnjfUJD
W8KzYLE9Wct+fr7HPJHAfaKHTkYbKQrb6RxBjAbE0ye2a4nBHStRMYKITJcQfIYMNxvj+CDLdsD1
AbVnoh1/5fyRW0U86ZrNC0YLMk3wuSNOH4xC7OWdRORJU5Crhen1cVXTpKKOXnTCjyo/kaKn37F/
lL30lX58ySUSGeXtevNGPufPdTel4Z9keLXgMgi33VaYZUCn4qpi4TiLdsW+ks0PNqgKzu0jbIoa
8NY8D/LjA5clxwBDss8ypPNsnwl3+k6OjoZWQ/EbjPboc3f0ou52tWPRKJYPn1bsY99WIk5cPJs/
1+It7m1E/UQiJ7XMxcg/ahDW/ihRfjUPyRYULjmfD7V1e95Xr2+ZJsgaD9odXZ8jgZsOH+eYaGqQ
9d/jjrCrZxjumWFJiTPps/tyoINipHIqgxAv+w9h00XfDBWD9p8ipjTglY6yUdJgOuxNnDWlAC/h
bLfBWTM99ORCnK9h8ZJdl/SxJ2Y50tgXDnRgBGCZ2TYI/HPeCANuH82nG8Mo/tOZKi97oEO++xyJ
34XI/+eDXFxTRREtJH9tixWC64wxd03tT/q6pSuwG3A0XfidOdeg0USiqG4vyhCKfHLzjxIeRF16
C4sRZUyy4jk/KIvdIziW+0nf+ot56hFZctTn0+GJoGQMp0Gou0giEukbtQbffSs4+Ga768keE1fY
3LCgiy6EJR89/5Gt5SnqY/uvovZpAWjFBrPmGFUqG9LYgUAHDNTA/urD0jEaFx6X9Rf+rkWa6cL3
aXS820NC1Tk1C9pyHONkw0RUUspciXBt7ftcFx7lwb6pkvKY3qA4tn0AGvLt5xyI0sfo76RvE9Tu
ha6SQqB1gfUep+oGDq/Jb9DI78IiesyGtVKxrK9YSqat+yxrX3zGFJIlvIEZzGAVApvbLXxD6BxY
OiZOgzkxcJ66dvfFq8wbOWsGumSyQGK+4YudPWYGy2VCyGsjteAo7mdnRS5Jp3pinm7MlK4GUUZZ
5mOTpJKLaOt8YLMkJOyBrEGhRyhBz/mCP/Of+oLtTguWETU3eGt4/zbT74fltyj76tsE6/HqCmJn
vrzusxMn+8MiyIcdg9xpyNFqJjvTQY3aTBQ2njVCoCshVpeC4R/cTiiE5L1cd8Yfp/mHxHVNLOGt
xEtNLN2T+Aqf7ef2vQSjTu9X6MPBpAt2xo/D95PmuhqOiXSUfpOaoz7cJcw3hy96Odz+ymDZ7eaC
7QV0d4nU4oRT8SmJX0epGZ3e5VzvKHGBoHrFWLUoGDZojuDVWjSfSZzxEVZeleH4ZOQWPWuAxQFE
15+p3Rok7o5LF/SEymf2D11kUlOauIHWf2Aa4TUnaHhDrLURvHuGtHiGdXoJMtq10aRGIqqxh2dM
NknbKXrqh/aqmpylMAScV4Wo/FydNjVIqmUZtipTKYusvG+8uht488KcpgeUOqNibtl1omgLiuLo
oQ/NdtViNZpTrnri1XE/mjZ1ctg8mF1DVpiR401ftSDQt5AHITTueGeMVhqZO/l+DKBdNB+ObFgC
gHFQNFTArjQJujt76QUwPyHsbmtSaaCcwHrwlT+qSdz6Ax5ibfKYWaCQCzZ1XOlrQPjxZIMSJqeA
n9U//S9mPptfcfTqanMaPlVrgt+moNEQ5atxORu9qps+uGGdhYKI1Xzm/Zzg+caeJ/EoM8z0AYK9
CiuVL+gObWMjzM1KnfYzNiA3QeXue1K08KZYvBl3c/F9Cs+jRGqhxcNZ5KX++YuYoOaqpf8F9JMi
gIzd0MxzH0j7wXz+21+JwVRnvFlrfmROEnI/NP7fK+kevqQclm2LwF9KdV7rHOZ1MennCtbFc8W7
bGWAc6TbR51DvpIVEaLzTapcZdCT/QOTwhTcYV+rFT1ZwILr+laXumpMB+i/jHZ/KHTMMqIvGieJ
SL8qA0xs9iO3fpOwa/ftIDINzEuN2Omgvh4g20+7RoPjeLuBS31Xpfi/9jhrIafUPqXHi6f0rGAF
Eyw4fNJy0a7miDmvxAEPHk+UXqPLB8L8UCviwq99pL4j6gOJTtIKSD8AGZX9aiBXb7rsY+/7kRS2
3AecQsDl5fbepL3IlbcEoHcuqQc04UxnZPzcpifqNWH65adudmy6USXImUJEAHAmpwo6/lvXQmng
u39igSdJqBNeQPBs87qxY9lOgBj/V8lxv4CiZpiDQxn7nYRagKW7p6pBSNxxCQHav3+wysctkj03
TZ58Gyw5YLt15wZuGjJx3Q8MMFecTFbJOtFuXA4wLOcl2k1uKgCRnbIZVXyo7NjQ7OOYPhZpOnvR
RYaqLzFaPGWmomoSFWki8BWOg3wqRYkaVhjmnEBrYBLzEAScrgSbdW8P4rYjRC+d9JHqRgyYV1eI
tV3w/o0g/LJyxj1vKuyC/mWztDqJOmd6LqNPa+M9wbqWTeu+K/FagbLCOYXtGiDJfDE0wVZKPHKt
Qd7HGCYCu/cEH2BL9XqfLQyoHs2L+EowIEOs6zEyH5pE7ARGvxoWuGBhL/D77AIimiBF1LbYw1T4
jQfotVwWa0D2eAIfEBLDwz2009duP5Jn2GgZ235M/yvcLq4uD1qOrU7aNwb2cKxy6MKp01UPe8I4
agqbmVQXp3kqSbI+e7Pz20byvprYsse6mxqcw68BcL8FWnPnI2vnK4tBG1RofFHJzolFZsc+M9NF
eqUKGHLveXti5PV6tl7LmLTuaTJswFSO9yw6g+IppEc2OI3jJZ75D+/fdnq8jIANYq4nawkQPkfj
cN4GM7clSCuwxB1ld5j+YUEWtGuZ2hDLKOTDpA3gi54bAgkGJX9M7s+5ypHJJxh3fsGNMaJR4M3H
Zxgr+UunVz4tz4+VIGP65op4NOICpU9z5KoGg8a6ZJMIEaDePhYtxH0hb1N/LnkkiP0ikewpq0lc
JmYfnfuXZDmvDCkUee50W/PNZ9C1fM2rWFrjC9CdQi2UNCHuoKlInaUd7chGKVObj3sV6+kAnA3m
T9MRtbsla61bGsQJfO/KtzgK1ccbmQu15Vh0sY17JpvNdXlJmiYxy2rK2pydSIyFdUBEzhx26M6x
hUtiCAzKFTIWM2zDF7MwYasgUpSZDZAqv3Ppulix9Wj8EjP6JT98ewd4GJjznxRqxVavleTOH/dU
2urVQC3XnPfnQKIKApdtHQXxyItAtfUgkZ+pWh/Zp2GivWstpCo045QOH6qLrAAhOIM4SmbE8t+Y
Pr5JgvuutbihTrn+W0R0RqtdrUnfCt0VFYdX7enkKBnJiO8WV144IjM0flWCdSV7C78GNttf6LE6
etFsF14O/hI22+8vDxAbJNc/H7xEmTKCWcdX+nJ9a2V+tzfTvAaog9mRSnSkxuMvXgfBvJSVZ4Cb
wIkJX8qUadEwKxyCx/1/YFT/KlmSrFWrptXAhdfGr4HVt6N/zaXtJ6XSu1us7T5D9nnaD5LTTN6s
9t4JKLV+RLqjiTYEutfOFaDc0ROoy/zrbXhyKDZzuQINOcgMtsWSWwInE4ec36MIj9HiWR4XNJmk
bBXixBCyJWUL9edLC4m//zlsv1ggTjct/jTvdDRn1+IuCNKOoynKPH9cAYq4b9jozXQGimor83Qs
LEtcbvBfAJy3B2qwr3zHygFFIbGSDwxw+ZAMroTl0le+xo0GzaHgAQAg8EWfeNDyzQeRiD8qM9Ji
ER5B25PuhpPFhwd1dziPjUn4vo/jDAzzcLwPJA1oEOgMLDespgU5Bf9Dlk+wetfR4T+79hbl96Fn
tJkxa3AXmEWGMNSQHcwWSLIjVqFQGn3aJAWpab2O0S1nlCY5tBTO21NPVyPbLKG2SD07DSrAggHH
RlOVYB0XqRYvnLQNqQAsqLOeuSKAabXWb8F8ZMT5q+nVnqcPYgfCxESvBJEVsTygBVGnfGGU381G
sB/Hf8D8uRaAGqoEjeSPBuivGpb9q0woVOpZz+L724vr2mzIJoDY33XsztK3FeiN09dl/Tcb4qR+
jAOgZI5LAg4dP67z2a0kbtUVd02lQasWUlD8O2YBzrhzaOyXX3VMQNFNm6DhCJA3ep4AMDcsBGX0
aaeuu/m7I+V/CRztv2rSHP/oQaW/Vj240Rf2G0iKEv7QKwsNAxpXMFRfVHyVXqPV2bIhUq954OJl
aXNDaNuLkgXE/G5TJmDMAoTMQkbu0c3dsjTGPBvfLxNAMSP3VDASDzNcLbrL6Mm41Kr644vdr7gY
uTi2pRlay06YR+cbnk08IZGRWUYgZloA49V5PsCEJTDC6ueTPmenngwkpEJnPMmX2LFwYEkNubxt
AaNlCru1wYgzp7LoE3I2uxkCHy9D+bsdpKwBfkBnqIClh3NqCwd+a0fZldeotgFJe5GE4H0DD1Wi
KOCCUEzA0yWntox8Cnc5XJ1llvovtX0YvF798CZoSO5KTz5NIYOp52sUCNme2Dj2D8+jqPim6HPC
Uge6I7sI2xclInEPYC5FrwjZLTCBbW5qqkriZUsxOq3OM8nWA2HybkyU/5RmE1Irpsmpknfyborp
hAejDyD9Q5XF0fP53vrX2DIBDjYoYJuitKjjtDbX7OGlYG7xr6Czk/uAeRkHVxVwNJmLB35g+LEl
chV7tLrY/akBdZWIJCYh2pyoFtLpVmynZZwq1WzOLrhd1r5YvEgB1Yl5Wd5aV0oy5DdacTyCRXAI
bzYCPQ+TKyGvUEW2fSJeqjYDdrKd9s6760ltd4jMhmfa4Jur1Rt4wcmGchYwpe458NdugNXhP2q1
nwAht81NXEIwbazJUNB2ehLjT3qrJHe019BDQQS0zGNXgxwBF7jcKs1D62BWKQ1vN8UzhitarA9e
oV1LIfowk+Nfky8E/be47qGUfh6R9phEAE/CmVlpRfEP+tK7AAsGhGLB5UomSK1u+cf8sEDhr83E
AFA/+ph4Je1cq3u6jlTZXoycXKesqv8ksk/U82rVFUnUCFCoE2i0eF5hf8lu/5Pa3ArwXPXf3SQc
CPzG+NjfqGCFiSoksnliq3m6qmAOstoPFk8Ec/zcmILSnjf9LYHwQfxKcpOmrnTMHorxoSG2wB4d
cfhh3GL9ywpx81eFDMVSdJTD5+vH+oKfoVm0z+gm60PsGid062vC54bC0A/oniSmKL7KFux3ekah
QEZ97xPrdVBM5tLkF8uTTjh4J+fIP2BGyDTLkgSSNpdw7d2WnSXR/wLpVo2XIdS/0N93vXyYqsAn
JGm/rvMTUzlWvXIs0dcoIllq2LR9sGziN65iGD0j2pnsHfieHj6aHPZUhzyHG47cqSU7MzFuSYFK
/h/e0Gqzq2rOvtBx3vhLSX8XTMAbd6Xs+cB5NXWkNkMqKFDC+N3rMel3uEz2A/R0L7Is8EsP1Jwh
jZQBzcVoINVaayzmpbt3XzIvHLu5d/v2oBvfWUcAM3WM5cWQjtZvA6kuVCshkuJyu1Lo65SnVGAZ
tSn/h4PpSnaEbQsr71qG954uiRqKcbFGSo6yVP4lz/MCChx+4B2A4+Pz/PIKcSl6smi22My+SsrM
g0KNd5dncZ6sbNwZ+UjGmywpUq2SLDukfTF21jiEc8tNul4UjQc+o2yUasf3jq6d+PawZHUc3eH4
A+QHgF8i1M3xyDG1SXxST3/DOujyYR8KgIpSfJmtteieEvMMiszXVAW8BTEEO0tKOLpM9e7OER2z
PvXKdlx2kn9E01XHSApTcZSsHlLU+xb+QFzOX7yRZhD7HLb3uXKa58lQDlt+vMhsdmsX6H1wgYDC
eU+q+TSgHBpe1CLTvEjRx+BwE1u86im9uTRim60kIcRBS0Hy2MoGJvSr3nlMgEa4YihLvH6ofQ+i
/k1HnSQTdj2Fh6XjnsGtrr4icIbWDWxJpQYQXnhqUteLAH/wWelRa5BFnLpf5IprhpXGtlTOFH3Z
dSW/MNe2N46fIxkXGTOQrdRrCuBp2aE1FRKairOr2BP8YrK2cLL6xmHYDAXvEhe3gfAPfxlZuW5S
kHQQwTPFVg1DHrumXchMduHF7HaTaINNsFPD/eQWm2R6dSNZYMPQCLipRYODN+2VV+ndqpE07g6G
Gyy7lv5BX6IiHfvhjrDQSHxhGCwadmgKpP4eFhHX5/eov1hQatbdWPS+xrs/MtFIFURhDxe/MrsQ
paSo+hFIJIk3x6NpzYMyXgO+mVM2M5GYGeDVcYDM/SbVFhyrYkFbyhnBffmjdZ9XO2ybQ+KNWd4/
P1TlIB1vxFnrnhKmSoYiC3jN/TqlybsZvxOd5f2ZdUJw05ULBDIjYVeOQx07UIpxgj5numKnjTW9
x2vEVbTr8hodkHbY3WAdy2kjmRAHrVGlMlUM1JwB3zpqH/TE1SgXkZOy6/FXqjK0OPOTx7lC9glz
C2jiYBWQhVnmuLmWqMPufPAS/vN92q8ss2SlIx1P0X7LSylzvPmcvpbTUObRwc0YEycKGK3T/szd
7UttHIfSyn846cplPFkxWney07qsqXt/TANmSZ5u3GPWdzDNyAJvRadwfk2m6wtlQDpmskBk2/zJ
9ovlV//LIec3n7qaUoLlCFxfnRCnP7kRNmadZ36kBvnCmzXBprd0TnSdjjnj0PagV3CtGBc0YhiH
L2Zzir+HyN2JYHd4tEJqkysKZmBDJ0ThCsQCy4KBjnHsAXtXptruBKhty/ucw9OHd33TcdQzFy0i
arFZaPmxqi/TmSELi+TjU9Dl3ET9LPkD5ev6xpGJmWgkUFqeK+hPcuY1731ie3YO797ugbEm+1QA
vVEhckUcLMPnSR6xExJ+Z9OGX7Z91eeslLbaj0gm1XkybvYf2Bov2xLeDZJU6PMyJDQnD/H+hloV
u2QtFHiH13vW0lwh+4MQf51KL5ztf71Qi2J6Avx87H+SG210/gMhuJSsVji7gSO9chP4WvTctEbO
8uLF215Et+U3j6kadIL2piHGQdv8DLU/OUm/+twDo2Nr2z1QC5dfg/y3aKAXSDW63/yaWaLNAQXG
UNdHinN6bI5IvpghjAP7S/VP960K3y1N/MRaxx1wA+M8K/E5F4UT21r1docJCK7d2/j8KJ1P6a3/
0zD05cdO8GgMZbI7EhEUA65WcvcjAPchdtiq/R+BQUlrKzWTBnjb/Znun06tfgXkJ/6iSzUfChxi
zVv1vbYWaIr6X1UZGtvTRkyRyquIRThp0CH/3LLIjXjKY+fS67QmVtFg8nY1VNwFPCpM9FjN132n
QCnnUMm197UkGcOfeHhH7kRl6NSpQGVeznP6j/Ly7mRCdiKUFXAi+KfROd12XqlJKskNAls5Sto4
C1O6Ss5GB+uh0+P82Pz9gSugQ4GfjQbXu2xQv8PpYiGKPT4STjlJBMENhAdJz6yjehYhZ4HIUjGG
1l7irIkvxoKQIACpS5F+HgT1OYtbouOEypNqshNBP0i+IMAEJwBvCe2mmfPV6h0aY0SJ2yd4C7Qx
IycpAOG+mlC8vIvl+aExJXh/7sjzbDBH6Be/sFkuEcShIhgwBpjgpw7l43PMp1gdnfx9+YVOZSbZ
8nrQ1JxcokPmulj7Ue/TwcZcPJvXwzBTqhpUcjZ5bL3lKiSpW0S8l5pYbhIlvhFh9TboSKBD/MpE
gvfhDT3slEqURCbxRWeYuC9U59UjZuT/hIHgNrCy1qtFE8v8xoQ8UYFfO4X3VdhlRK0C/fZger2z
CCxYK4+ZPXkMSdnN6s8WFPiWRm4tQVscazeXhcryJEGO5yEkfLtVe6MHIyI8zui7f144Tn3OCaDo
YHH40ooeBDqhEMHJGB7YlujIKwqw+CVGqHoCX1YmcISrXdfDU93bQd1ZOQzz8NreX272KJWS55pF
fOHuPAGGUZHuGECoD7MjCE+D8H0y4VyOhqon1BdgZtqp0mnZcPWE8cSdnDd5DSmEj7TnlzIrASTW
ktkz4XfZ7PEuNmRM+WGyx/BF8Ba4isc0Guz/5jHOjtAlfdeS9RuXVIL37ttzqOFGGVcbjlceGsrV
VtFPKe+lAiokbE1icd4l48o+vKLSCMYv9WopXrFOfm09OjutWtsE3CTFt+7Dxws8KsJV1MJAQymQ
MBxvYvkKgr8iNWeXVABCJtBjI3HGsFcUxKCYtgpEdO+oa7lUHObbW70YeMkrCj83Qifm/AIOiykW
v4DhKgFfvXbU1vw19sQQN6NEfNqaJrdVKmC3+BbVGmcQSqmRDNVwGnl3oz8Ww04irr0WFaTpYy7T
eBrER+3EraeTxwMibd+VMAGhIpfPECJ7n+evvUNgzaWy3Cqy3elP00mtAWcyzMbxvUncjKleZW2g
FuCMC973VSYLHZO/QOlg6Cgw8ZJq8ktvkydE7ek25ErQdHuFRsAl273OKWurM4PAuACmycAGpVaT
4rhNr9OLdw7P4004qJ4FenNVsofGuJmwHH7gfA6K/FeHVNwqLKpyzmzyY+Map0W1LHLwQQDbtj7j
y05gZbSQ6vy7hlz1Oim4MA55oNuxvAwwRK6FSqexuo0QIHxe5wR7gO1EqOxlZ5071lFHiGtrzmp+
uBo7VXq4sTqyBkjGGKwmmrz3NvPP3JmwFEIbqczNh6BIBluWsME0JpcG8M7rhMNjcv3G7Tlw9S2J
M2DZXL2j0SnAyLOkvKa2Q35fh+JbDvd7zJDyjr5KWZAlWrKeFfAPm4Mi1QsgfGw05bWUMQqCw8rT
vycocgjIPdOg8bZIsNGN6qYpa2W0Uq26Q264vAI/0X5qyRBn9FGtkZKYQ8ONBYf77yaF3vLDKony
vSUHs0NCBwo31CCSfkxr5Q+k7GDi4vfrgSDJePUEjVTPHT7aNr+nvhfmMcyLJpb++PwiuQU1ABb1
caW8n9h6DgGIuhWxegE43hDP15pGC8v6suA7zmr9JWGxGYrpTrRepSfWsYViaotkOtLZpa65Xg0d
BQvapdaHeaUjiwmgUer/hosxaDqKo+wVEWIrhLJp+0rWkak0Wdeeq6Q9zJAwiWcgu8VQ+sTTbWfO
bjtXSHS94yWtROlo7oKGTedG9KvODtUWi1p7BhqyQSkdfvK6zmA9a9GLNeXKdA5bvzJb1LSOJAOa
7ozzWTA664z+d1Wv/unNmn8TCaMGFlST7pS9ZsNRu4H2ded78sJjCwxQ2TCWoNDe8cP6hId7WPey
3fhnRb8mH9hyQS6tuvgwlyBYW+y/vd+Y17JicmhNwA29PdXCaZWl0VvTIzFcG3IEJwAqEhXv4wkg
WiLmbISyGOQ6s9S2l1aam9Lc9dJ7ipeVgiRTV7cuMQL4fXsXRqsJpeD7pf6MDFid3aOUY8gb28Rj
OgKODRdkDBBHQ1YidEMnKA3lmOXsWyQaG+QxgpoXwytMdNbqS1KGlV645yUfbo8pxMR/P66X/SlR
Q1oMq0k0MBirjqHXjsJsZFDyiskvE9DDKd7Mej4BkwKM9dilBEiHHSG5Vrc4uE0kTDbVE6Jx64Td
qfs5XaFoX4tusR1ZL0DgiZm0Cyn0OtFCU1iwwwtA4xzEsUvvX/YuSmGxOh7JUVbkW8ERKevvrLaO
YTc3j21oMq/CO0cSvc/JKiA2JuS44eXkH8VNveDQazsJQ3dw4NC/VfbRKNIxvMDM5oZGN3+HF0/5
WGZsugILD1xglAmBU3WCWCqOb6PFqKpZqKLsMsr1PHnkNwNhrrg+K4aQQ/jNj3SQAeU3CuLQkxms
MLiiZmEcqUoCb6CCwvoKRF+8lywYwMfhDzYfOv3t7mkBl3DpdU1egJKz92oByTIy8rktv4BQ+F3s
tYCxAQic5kdoGv6A/QTiFslEVG9lXISb7zLgFWZ4BW3bLFTtPDts6YTp06504Omn1Wtn3i5ENTbW
evESrgkqfBHqByYO/dww2C7v6yGXIiEVPFIHxQhsA+CpTjRcTBscdsYHCcg/2bjk+tiwhSdaQ2F5
xT2peuRAC5BS/i1cqvymskpXRH5OFBYt4yTI1aUYB+svL6xw/MwGdqTJWJtdIzcWFwRCJ2Clgs31
V38ziZUOtNCLVlOnfen9cyfp8tWFtmdrEEXvQNnMScAL6Ox5bJbwaTR4LSBA3jHgfsHN7Iy5TSS8
50xiSpyG+uRvmbi7AXsXT+SMVBTbaZo8FNjOcuk0dZ6kWNUhbOQw1rD/WkuHcvkZIskQzWHjz8J6
DkbLHfFT13Ybpref8a19x/ZxUgWXpDB5ZII4NjkUq1hC5mJCgC85ntCBZqYbCuP0atz5mtI4Vdaa
fA865x7QaddnMhAW1+Xmptq83jgrwwqwxZ40SPBy3UjYkKcF12Mp6k3IgtRdH8jo789JP0pxcjcY
LP36n5CuIZqtKc06In9p7+cbpe5hYOGmadXLDY3yAulZiQ+4PpiASPrumWO4BhgonCzq7c3J50u7
w1xovXpFP+wwTaNxHFsmYtZmXOIwBtGM+6geyrRmZduWOo+wX2Y+AtUzcbNdwIMPagN6s82smyaT
Nle+8h4sbWN7TmWfiWjept5oVGnZugiI2ddtxmVi44Xy3Oew1eAj4V4mC8CwvXa7CXRNUw/7LbBw
VYY9EoFAItmxIUJKjWq3dP3s41jE6b021y86scQqSGh/ap3R2rnNvYjyFN8Zje9k7+AsN3gVAqay
LZBrUE9ilxY7QJb+8LBQlm5DfUX1Yt2exIcTuGFhCh8OOkL/csDAq7AOvnmD8ksMRfZuftsqouww
UV2WdcBVWn7FuOcLDZzLEMKahZJx+XQsg/AIueTivaRzNk/xn2m54WFqw3zNCRuQ+XtEnIEVr/dA
VJctoX5RmbjjdjvY7YlG4j5fj2jkjPUd98mr+VFXUwhg4351WMj6Bu4mYIqBQh0VtXbGF+6axrr0
jyP0WybyB2LJ1YqwFx3cWfUz4+cEdaw3WGIPfMXAIWcG6OqV0g/WAEp4nkVrVi89sQaJW5g++BH4
rvzeaKIvgFV4Dninj9fC4/b+g8RUHzHBWI5GN6GRMp/KJP6YsQT+jnh1KRn0hA4W50inTdDa9OqH
xpdUPKCJcM6Gh1HW9SIy5HAMu+glCOWhlFojVkTflbaq9sBhVsDCUtEkq4+zYWb1sUZuH/SKvblj
Yg3tKV9F0opZ+u0HUi4nNFieIYrH8/6h99r90KUPx9GI48QAflEP3SqVFFAcGhG+Cgz+isP1AX0x
jEn9zAocGTgfKenx0CqljVOCNENACHYMVxzqMha050CpUtEQTNw8x4Rs3us6nhgC1UMaPim+spt+
6ZHCr0/4tZBx70PSzIgsQ2/188vkFl1sQc9b87cUpcm+PaMdAWuDBrpnSivgEYzX+vx5cKun9i6s
umYnsNLNQ1zFGmBFqQDwfm0nh5DcsR6ofHlM7W/nnsknDCURnlp0Vi0nalPzpqmMPeL0Nzgb4GJz
nyuGwEmukF8NBZxUGPyeiGkUvPOly+5Jp63rTeueUCEjoWoKTxmsHudGqsea0SsVPEC4dxvsV+xF
+Dy4x2tD4SvC6EPZyXP0BBdacQ9CwgFqqk6MnhaDjmYdn4WCEsCyVK0SNMzXdB5WvZ/ynuB3Iy0c
u23Kp/Ko8ZZa26WbmR/OPrx4Jm3p0FzIY0R6qtIDdYHT7XBA9pDdis2IMHC+0rMO8G7m97cpXFQU
mKLcK7lTC4qVZvNYIhRjtZZj9Q7cFoUaZCIQFG1XzljZRfogCPQ/2zXh2hemlLy2uSCrTkRXI+WU
s1X7dldWf/6smhXUIXZaHK6SwrOGyROyTf7U1ZQk5GJgWyQ53pI6dmdg7z7+U9e1Mg3cgXiU6yvt
7XgSM1wo98l07/QTfGGwlJtjEbzbz/70NCXaFJf2LOXWqAttF3iK04jxoXKT0RJv9GUe3mNHpfje
lkjRNQB1MfAgBBbak3sMCsrjtRdeVujszpWwyBnC3VnYJQqB+33IqymB89XapUu8r+XFoXPA8M/g
EEwUUO+AC5TCkRCmeS2yxnnB2U5jrRHIFeJr3D6xtxCrT+9oUa/98NqeA+0uuGGIH6Tnpblgis16
fj/vYkBDhRHR9K8oQQ+RCcxHe2PUBXbHbw2forPItNqx4tx6Rd29+7/vvBYOpQxRR9lR4pAzI69B
GG/dtRmxwOfEM0SOQayIs9SYdCCffaMpXnLKvRW+pizCx+2EHRY6Mrx4L98JapRKkzwT4BJFBmT3
vVpoZHChBkzw468zKO1cOtigxPLSKlyFLn0HTe2U26UevtLDWNyT13D14OqfDXjmZ3JoJGGDCpc5
v1X2pwS1KNqSIrYj0TAanJK/DN5C7lLUsZF6XQig5XJDwZ4Vic07y1doPSbFRZDogheAoMcOYMZm
FEY0QM74mMTebWMTQObtvkahMeb4qEuGES6wcVoH6mMiCsGX/UDZAv5iLSKvR2FKGo6IpnmLSEi7
zf62H3gbWp+YQFgXGlhXIBZwbA8NX4mGzVrc14dSrbqL6AUY5DDtq4MouKyYhmqnZxLw2jPAnfgE
CIGXWphr07WCsoHpxuLdUc3DFy+kK9LnSwymut188JNtru2s5XN8tM4eVwIdkb9DmXV6hkKu/tU0
krJ/jTxMznWbjJFfkbverkQKv+QbMZyCi8LeCA6PSaemlsaL0yUa0nV9meRFwC5iP6qZe5k0IVyH
iAzR8/vPHSbozBz0HV62hkmjx9eSaiZjYaBuH+gDxE5PFqt9nbsYMBZHNpdi4/gzQEX+WrqE1SlZ
+NKqUoCfeAhBF1Qk4Vysa5LVtrwJGDYb/i2wo5j+NFIM6TWtwQiDFLGj8fJyJ6Wce8ZIRfbX7hvy
ECpN4eal/HyK54XxHgQWWb+NTRr0yUtG2jS0DgUwHU9DUTqSzQBY1pT80hMaziwAPFzmd0Ad2kC0
8jgYrSv3Vj1yVwFzkasTksbfwRUVzK8QCkXp0/P3msLmDyx0hwljKtPt4pYpyNWmM1uPmR82S3+P
bbDEcILyjV2DDAMVN+gCbL9geLs5Ci9+NGqNQ9sZ/cjmxE8kmBaLxYXRbwvPkjojTElmSyBfZ1vn
RNwqAOeTobscRPN/ZDZJBuFC+x/hTK9nacq4U4iQJLHOV+FCeZhBuLFD+6gWZVoWOqh84bvDBijq
38G4h1XOh4Cfzr+Qf61tESwBJgBVuYIGmZwcx5ERGshPewzEHuhAkZXqxrgCW8dDdkauKJfkN2bd
zEXnOz001Eu5B9a/fZX+73yST7d29hU8OJmHjD2J/n1NUtHy60LrTE2RoL8yOUS7+SUrZ6lYntlq
g8R3cWhgGPIi5cMuUsBVHBTzL+VkHLwYgU6F4h5XgXFgQVlwCnEwi2eImNbiBhdPAC4bKDgsXnjD
sAmSY7HS/9atjsmn8fWx6jRvO4632PdepG+fvsXfD7wkG/DDBhrknYmntZMZKMHilnSJpk9Pqk0V
1yjR/wkOBekRu3Zi4Fm1CDLijwnO1c8K97OzMLTEJjqVKcqgPuG8KLQiR1cZTINzcA/0ztNiIjoY
rEmBVGnbHEsC9EHg5jj2U3umm0Ge/trfaG2pvziUddumGwr8cWi5OyuD8WYCnio3capGHwfJUAel
/xiH8GeRWhgq1VEdNTrvSxO76kBCHh92OLNs+LH3DoJZi7hmrhXjADwswC9OxTV5/qb0L0po/KIC
HobWHgae8VmLinUffdiwA1vyHNQZOPEkWH/ZEa4YWS0UJhX+zzFWcHI3zm8zg8Hyx+WqYWGxBEQI
qSBP2Z8EDMSDBr1iM/dMsLMf07j4IZrU4+qHTLjeg/ZXqoZmgeTFLbLr0clFEbhwMcKRMR8cPO7Y
8v2GJMrEMymPXsQFcmxqiryk7mw44hkMvFq6plzGlNiaKk46R9O2uxhHct9QD5FTYlOr6cPR7UBf
/ar+gKyLYhpdn76+ktD4ZnYp5NegVP+2bQ3fsl4kpb5jCGMKLOhcZ6j2VUSKoxZbUnRqH7IGU90t
xzRHAfqJUShbJVV5eQUUBLhMP9DBWEqdH7EdDmBw/+wd2kP2a5DC6AdtLbsB/PvkB7sIh1zy5Kok
LVBCzTsdfUdXfU3zDOAuHbOVbJBeXpCLmPzGm8yz5TyOAbUJDf633PetVEmbE0Vh8ULZWucpNI6X
G38vZuksVVrH9IUDItCNDPBgMrAXx/rxLns7I+CZv2hFXyzr36cKS9PHTimIFqZ8x7zMUlm7kaZx
M4bf+ol5nhxn61KCrTBZ2gfV/2EhoTB01aoMvFyrkLFp8SZeitLVdmI264r/Y27LGzfvGQlb18W0
UNY0u2OHvEG6X9U/cpFrc/gCXYNhK+tJm51y2paA+rBfw7PqD2VUS55jxyWyEt3PycW4duq1q1tg
Sv6BJD8VZ5Z2IAzGw/csCLsCc9WPvj87HN4yauBSzrZBvHjPZHP+e4Kq85KH5tWRXYqLSCckU0QS
ChVzr2F7r1GC4OyQ6W3nLxcuYWVT6m9TPBtyUHSBahDYRtQTmZ49XavFEXujVKTAR7vAyZiZM48r
mI1i4GRUVBaRCawQeIWAYZEMRMHA0dxRnUqgXaCD5Jh0OWn7YLemRVfcr86C/nlkzHn5dfKCF5CW
i4hAHjzLeFTBwMynDk7RN7pLQaL0TupBkzDRlncJX3JuQORSNeEky/FiPBr3udRLFndQSTzDnbqY
zZHe7FaJUOyj/8Vy8Suyz09I/KyCVmc3oIxqM2lr9hsBKgZGPi/qrBhOaOcIPM9iHTArNomg6YAj
MrY9TlKfgQYsSucVICGh8kCXN1qGUGREwysIhD698YWF11Ifk4c/AOIS73JYxGaDTKn4XS58L1Uf
2bH7yuXfb3a3TsvlIF69sk8jN6ZkJg1z0ORNWPy+Rbg1jS6idtRh4a6sh9w/1Ne8wkhNXa5F9vgM
CJNIwsEzlAoD4WYBe3Qr0LxpIPVGlx0akEdoSdeBT0Tre2gEcYmzurYqWgavHpoiLwJC9t+gLwE1
ym28fzwn6yNKqOiYSPabSai2gXUDnUo044xdRJoRnfpDXcPNQsIFCwv8Fvx0O12lPorkCSMVMmOk
Fyo3TPmR4DuIrVNP/8nuqDwi7fR25uTgnE91ldJW/vMUQQ7/VU4cWus5vV6EKfS2KZ9c4oNX1tfs
+TNKcR7w4rNymOrzfnh99YRLvCNNMUNXaiadFq4+YweRh546mfT/vG2QoBht78T8acYXJj+QaXuR
XM3wIVFvQcKjeUvPVfBUOVZo9Ra9ztmgN5L8hyc4mYsZOHrFiUws/VfcGyCZg7YiVBanf0f88Pnb
FUZkmHCZNJwVVsJgZWW7KNYOMljtrQ3J9aQfc/TUP4hFSS7Wkf3r5Ws6F+gAtp4SIzeqTJKHaq5L
dsPe7ho4qobGtT6X1i1CAmzJmirMQlEWT8Dghu7ZZnHgrqHQMKtsETHAXbPMjxyDg59gmZEdXxVW
TMh2eh9TnALa6MPDsppMouYVR/OubfE4ZGkfvE26YT2lM2r8wM9/TpClPlG9XSvNqCfla6Yizola
G6eiDXFgfVKAfWg9/szWsAW68zXS5Yuc5GOJn+G1SAWgeqtch79btLy3SBWpSb77Z1dSDmT+8l8o
5E8vFC+rnmDjINDukuT+Ghvs1bapBE2PvWIHnM7zoZ84HkVVl2Jax19jbg3p1ILQZ6s3uKD2+qjy
BQWWkzlgeIjFjftm/xVwJcPnC4NhDo66Xctk0bBhvC51bx/rv/MFFARbyXYr6WeaXN63ELEmBC0G
S7MTl3h74b/JOjqp4/cZZOkoWbpvGzSR9oatHImKQa6FVWcxScPs6/EDEFT+pe/Wlxpc118QJjI/
QfzxNnNCEnE/GE8nmwxwtk16HjLBfpfVo5HlpOqNeHd8hq/EStYjlsP/1KZ9v07GVYNUKi5NXUpT
tN+53KXXvOe8bktRtn0zoeO11t6zxKS+5J8Msu7td1KRzUc2/U6cOJOSkge50tSzDkU/JySdQuu/
IzFqejIVrDHU7SRQHTBDuhD4hb9wvd5acSYvtYOd9oCxAqcBrt5zKpJA35TgT3zbo9bmlEFIaqnK
5vz0V1R51cx5HGgLDc+slI7zXL9IYKoYk9aUbBKwx7hmMCyQxhfl1iFG8WHblNTMYEnLGjIm2QRP
aD5Bkpzo4ct6qYsWtuvPDigiY2OlHnrEVOVzXbqF5T5jBgbMicFZZ/vH9k0sdCVFzfaikKmpNDbJ
mwDFL7MaM5X0v4be+51VGMXJN/S1SJ3PE3R4AHmv8OWFinQskxf6DcJ7EpsykfOpDAwCTA7D8gsD
CJmFCwnlkcKeF/HmnoQj5KZKjfH7de9usP6tlGAir8vtwOG2FiTDiGC9HRBN3sivK+gFaU79KbZu
Rv9DA71lVl8noPbc2zHK1TeEigOHz5kiREwPOyRWyTbN4VJrniJaay1b9NQWzMVqKqDBWS4/fd9g
MyS2PBXPb7izXvdlQfBbV64PltVZE5c/fgi4/8WGltHFOdbztr3uLstmcCOx2YgNF9wnkG4m/cVL
mSKav/SZcwwWf1JXrhHmMGAgu+/q3kVirgIP4uIYU9vFCstwi1M7U1ZYMJk2tGAsgmT1/l0XaQHz
USCXHhmoWlXnRpVItNt+/q7cnrkUy2yh0/0T+q/tZ/2yMvGcC8JwckH1inswTVrBeTTJVO6xtSFF
aZ1wMWw8e06uoqW80/rB4LBPfM79w4nlfXEDDR95jKGUFwFrGDwEEk/W+eKHD07lM0FITuQZrYG7
JtzU4oK6FcRGjZAFeFPEaKTH1L1EcU/XSyZb1e4mWKcsbSW6Br5hTFyEcxbWFY1V/qawH07CQat6
QTAzMzRg9lVgdjjmzdNJ7UUOpS/YHhRWn+Wlqf9qCWICMq2iNzPVlSmBuHaBEKNzWRHskxA2MYTb
iX/ttjwip7QBXmLVNCPaa9ij80KUyvFAhAUZ00lyRTmBUf6wSlJOreVJzOFvfMFzyanKabytsx5d
2ZNQ4YfylXQuGixjcKzo9RzEekCCktT5PH6P5lPsit/yMl4jbt/IQNFKJh2nbZqsqezuEqjmbNpf
RZ9TQq2PnD4J97eXSMy1roVP1Q7YhLjk9YeXo1qc8jLKmYpE4CjaHz4GvYNLC/Isgd8mzfCejCXg
3Tf2jOI00+JpWuVqbRt/DsgiNbd/S2v23leHpKaPKMYvd+uIAawN8Fh1l+LGnrwZWClIVx2v0HBy
mL3avtu18kRXJI/nks3rs6IX9B6kg0rD5PA5qxErgP8/tHYCjJA8GqhvW5vEsxpNSwuHor7zsruE
jVVYvRgRdGqGdvH2n/LFftLjoBj0N8ca9BYISc+hcd7zymVsGZp0ckjEAhSlLKjHCmJOsObPYlip
ZSIee3tbsi/IO0F79LV4Csru5ojwmaeIzyARFtIo2BwI9HKjHkgnmTw1407VOA8Fv738W6voW7gO
fZbl4xZxx+KydO9ZT1Wka4yZ4FvqGTEj+i27YItg5FKIs3erl1CRVbbBVdIDPx6BGiPpytHB6AkJ
IB2hdXgcUs0/f4xwlkBq9oMLA5rHeRcL/EnBbJ59xDWlYlVTaYHkJ5PWZrBeT9QZy/jdC5MQngKi
cBsMyJmIF9pnPhgz3J81AJqoLESn/5eSUzTpehKA3m6V/HzOJe1WXNgseGY/GxRVVt7/Ol15ei2y
le5TPw1SG1O5VUn3J/LE4IX0VkZnMUC+S30UgR+ZX6sP5sjzhL/nTL6xN8Se8KIplGziRt46c97Y
pVKa6S3TdrZxOSvAhKQTtLImp+UIhq+9lNEti17LDryq7tYxTLX5PE4E4hV/KjVuHqH7YA6KfDni
TkpqExcFP4VKwOdrSNJDHvqd7ujQBvlFhrjelqHjhktdgvandJFBC4ZjXvd8j01EhbNgZAZoj0Uw
LWRZYtc0D26TmuSU2y2OF76fnfW944BUQIsWN+KA9sXknkZMXjSiVNkmpmSec49fh2eFCv6Q2UC5
XC6Mq7nkVTwgrAvYiFO6xs9fOmJya0XVDkBzHwXg/onFmEbWboWlIeSZVhcra/c6Q2pdofQIiQLh
3HQ7PDwA+2LKSPZsNBetpsC//7ODsaRVvSej2/Ywz4Q6BTeH8jSKZVM+7RsDSdY2O4PngIoPFsQP
+RAnjSWG6AdJOqoykX5p2OEzQ/AlOlanbG2oaishW06Lg0pyxxJu3okVwc22Ju0qg66JrgtKpH0z
Onexj5tiqj0HCNvpdMrsbjZKffGYf7iVsDUuSYIcyab6IVHadi+uIWh1hpno3MRJiE4Pv4xqiLQd
66Jp36jHv5hC7orA3yo6PRLySNeqJNQBl2JzLm3WSRZEUf7vevs5u3jeIKBrrPIm/7yFlQI3mdJ3
jUyK36grtEXRdxFWLfLzF51tKNUAZjolWaEQNCx15ZvB21DiN2QvDqwUY40A1ohE+/KEqaShrkSO
S8zxtHts2UpO0C1LDqrxZ7vhJ0Q/k7eKhnyc4Um8PwNNLx/dCuGsAXCuTArheHKOh1BTy4guthDv
xlhpblkxicK7SI9S2k0xn8qCNatILslg7JvVJKYLzxBvFgSUUvuydnHpq04msT0SvWqYQb8oLMtj
6pM2STf1IfhDihnKfKnJvMO8lnWhMagvdmtNZVRhdzFzr0nZ3TME0oZp7He5qdf1D+fc3dSUm+qG
tDhxDtxOMCRw5lFw1yQJEpGIHpUoEBNIHI7VmUC0rg1ROQWKYVlBYmsZBYxOjJMbxUdRmwbg0uVU
bBKi+VAAz8uOfnjqQckJHlViFUgvzjey2FFTYOzU7p6FX6l9WCv5d1tFSfdoQ3rV0BtO10cc0OVJ
Z2eJxxKJqQrEcemHbB2e116jVt7VuQFpk32vRQcR10bF7q5AEWvn3S8elCTLWUdvJUxVkHDAflaM
i7A+cQaJHEsC9e8TkAiIw4Hhz3LHK3REb9R+EeFOj4O63mbTHirptDtnb5zhQcsELwLuqSeIVkDK
FAlVs1ENwVgVERkS88VBx/ZX/Dxzz2JX5jMHC+fU+C6SGJGbCQoIodEdCnspqaOhPsQuUsVJzReW
YiOkzVucxwB3RQUApRvsWCUHsRHZRbAatkr5S+WRetU5SMSG1FnlWmNP7uIZKQ0zutLMUFkbLGDD
dVY/l59z+JhXkI9ajWdTI7HTm8nAm6mVeKM1VGH6U5J6fTwzPeJdMFX6OFN5A9tC2PJZ1Pif/a4O
XZLnYnwWKwBM6ke+oMDQKkqxMWI9ecilPKr6Czbojje4eusqZE1oignY4Ic9zGuZY320AqkflZEp
/cjXfw8GwwQg7ULK7/v1hAT/ZyZcoLa2QLA9KCzUHjamaeJChyQiJmfx8g+S511VSBw0Gh56S1Ob
85qak8Ccl6ulGQUAxsBGdJ4M5YrAzPJ0PJkSbPIanY9ldF60hpaFsVBhcxTwLKvKfFY2Jgt8g4fl
BeHzAFB5UbQ60YZKg6x9cXxIS2GDOIr7K9/znqWAJGynQDgyniTcgKnHdDgwpqEMt3uUroe6KxJj
IuwUG9JpLiRfWrQ5v6OIbVwwSu3VSJsU/3xyng8eAb2QQ12hBQKkK9OXJW5ErCn4Xt+TeOzrS7tr
MMmA2C82oetA3LOBGpBRl0icycs84BX6uvCW2gRp8BJaF21yFmgZML9Tdb/fmLYS9BQ26DiBNnmH
wKC4fOOL9uihPn0THzwCNICZqmab3fL6JVnZamh0E8Ji/6L4mqEkth4AucC3NayKvKSb7JlHqC8E
XIRBCY7KP/NpvOiMTnZVyxHISg/L28ecfMXZs5S9RW9/7uwMuX0+GCcVzZU1NAtkdLRcbfeBxnTJ
pFgXc7Cm1ONzvzLp3liicz8jBQcA2XwE0QNhbW9yCfzAYNGUCp/CbkLvSx3F/toUXhbZKIfr9Lz7
fFMweo34KKsoOAmbYbu+5tAGTPYj72cLJmZmxxOKDyWPyFYr+5rTGTzZzY3Yeb8epAemZQfSyzZ4
7VkG7kqnjvfQroo2P98/Nt7pQ5Uak+UA5W1qB+upUU0Tf21ZwpUF41v4bt1BeF+iLsZX9BXL31Ym
Co9S72yZEZYKBt+JD1EQzCYcSMZJJqPWOVlK7G3YDy2drWdoBIuysiWXRrr1YZqfWt7O4FyDr757
55n/NsxxOUc5bLIsWUmRW+4P30vxnbq2v8G0y8COJeeZgO1XaRZnPVUd4KT6rSOxKybe4ba35r/f
FL7l+Ij1pM9cUgSMXWHCzFjSeN1zJ0q9n+UVfn9UhzMGyiAMTMmMBh+CElTFqD5ndVSlTqgVOJN0
mswi4S3vdf1clu/Yz1k6pMD+/vRoqakpZhVSWaVYjmPdpKGZMTRQWwhNdyN5IrGnoZrJ7qFZ9U1J
BzHju95jsaYVLCQYoGNjHwpP7q97kSkHrIPAQuwOB+c1ygLu/IzunbnUWnZwjibErnHY2eYAU7VV
VjnjGvpWT7XcShwIw/ZpAhvk1SObjyIQA3knZ9iuQYs4ZNug5qN8bET9IV+Oy7i1dEoEoQf2Ajo0
RWJgx+QO3X4lJztbJJ5TRWJ8mSleeFv2NXGt/xfevcXVIs8fgL+xPwyDSYLhUKh6z+hKf1XcnRzH
OzAD1PrB/JVW7O/lgGPMc77jVa6Myy7orWZsM9C8iBfS21d4xhuHuq+CDbqnSs2YXhyHj+h6bQ79
AlZTSt/+8fKhOwHr3nLkCRkzOt+F+Ykz9AIv7sPdQ69fYPxYrsbhKikq3a7RKGQRn4EdE41xa+Iy
9cBDuAsW8+pF3uwE6L9xVkaOGOOV0tWYWn8OaRiMnFjAC7XLvRpfQ3AT0Gj913OGBI2gA+AGlBAy
8XOGdNFgRw6wk6BJ06NQcL8FtPPV/zFqpDniKT2XsjhrhDkYKvp4a2Og5kfMqNx5rOA12QbVloMV
SHpvNQBtouuEm/jnKhHjhpAmJTuF1bb0LppLDCwRSvFIZYVqRKSqkzZ0Wu22cg+ln0XWCiCNMAz/
naDDPkfHR9dDbT6J63y6camGbTHaF7DsYWWbnHK140NXsCvCgyCddnFEPOjhPZcvBL67C4WvIVsq
yotyUUe6QvEFL15Fo5+sqZ/HqnujmatqcWDuMXAIGdwCPNO7HqhykMWkoZJUd9p34/EdKEAELAa7
AHjjPznpdJ0jd3cNZjS3PAbUFE7UzyNYtsfWpHEsCgc1huugmI5VKYWGb+pmKToA79y/sxup65Ru
XBoatzBuJOM9X+bvu9r0MgMgaela6kKpIisu8s1jYBiAqjCHqqkDaRMRY23LJzw4JdLrl5QoHKBi
5oIZfHEHEoVr3ImvwBweYjvVxjh0ZoLhLjHuBEsugkrd0dKCHkq4AKiSdu50rPbIBX/20Y0rzc/s
+yhFHAnrFIDYvS+fLSggd74ukDV5whDqfh6b+hntEowe+leg2WF96oCvkKFM+K4eN/HwOMaOzaSa
fVewJhiNWiTyneqT8+nyCebej8SCYkG730YxAlUvRTGEAMDY10MLkAChkNFtqaYNl+V1IV7ofxzX
YFgWEED637U6u4R0pLZzMhFPXylWAHfDj2CMmNwmOjVvfZMMWmXOs//B3BdTjpoDRijoKbEWQNUj
36YILNwUMNby/APdAFVUdrPuygpuHUY3YlRyXmUNiqgFsGeBkwOlA/M+NBd08toOOpqzu3NlOnq/
F6uwjLhlxRJKcb6fv7+Ee9FPhA5ffLuAFn+a5HZH8dTFOXzEZmwGzqfr4EocHovIDwFR3e+wh2xH
f10FDCtK/wAUKsp1PdaN6F4Ow8vL70XCTHayUmt9ZHMJN9VX/PCPUFpfcODFl+CMLPRV74a8nf4R
4KGPBPHRQbFy0sONmfjulT3bUx5k9YtjiWw/J68l6SKSbca72kdP6pvfXDtHY9PnN15q7i8abJj0
SC3OhpTurIxmPVn6eeaybpLzm/uLc0M2W7Ux4heVPQbQhe7lJ/kfMXLXuBuy6qS65yhZ/9VlPolF
ksdRcJzLvQLma0npQuTYt+JThMdjn/Jx9L9yg7QsJlMcezHEc1S9jzjezM+gqYTIOHXmt5k2XYzr
X/4bxUFvM/kzVnKnTxlqEamLniFiWIkRxcmWdYpBtNx8QogA6qitdwVBt+4iUF6HGkp0/azqhjj8
wbR2UfHSGAcWMekiewbGu2w0XmVEQc5H8zFqUzkrSzoDHWj739ASPWrhtrfOSAY8Yr2VroSSP9ZK
UwjOWvbvZlO44vNSToW+7UaWwzbVlrl0g99Kw5XYO4pJbWTatiFJfeoyjRh571QwZ5PSGDGtAsgu
vuuYw9+fUwavybPBIno4K3DcnF+QlAUba3GF8G+3vgrXlMRNYfJOf0pb60kQwgSGV2XNR+C8f3T+
bhrHVcS1c9z4wR3tv6/su095PQ+yQJeDIkDalGFturmic5oBjtw+N8wEADUP8l8Q8zj0F2IMEKzc
QrZoBc3yNmkDZaMDtjLbIWOTZuRoent6KFrJeWyQpDbsKewQJmb/pvRddSR+16iwTQLR+k47Aaie
2x2PD5n6NoDRyE0z+SLcRZVl5RPKm82uPLKZSP47D592P2xN6OnCMnkamR4nZuOzfDXtlBpsVonN
Fz4sa5j3w8KjX3kw+ppyf+/eswW2IW+eRf59q4LGZJLq1+mFgDAaAEQo8NZtSal1VgBbOC+wFb44
/lNfj9UHsJMC0gijLv3Nr4p01B49CUALbPwLVn1mdgkaL75HgpSqOjPFYj3PkfSa2dBt8zS2CGGm
Ofed1sIl/7RQ7YbRnMmeVzsMUYKsOenvEcWgji8BM8QnB3UI3GQfYuOKo43yHIHV9PC9LwOkEfcj
DMwZOK1Tg/ijCWm7zpXYUFtEVI5o391SHkH74cRRdJ1ErB7akt3tjkM/wPczuhiIJH9yN+SNEVZ3
xMspmVMVRTdhFcywGwI4k9/7Bqvyd1ufis0Su42M/21lCOg3pEWaQQEss9fkfnIJ5MRh1/3yVMOJ
IWwVIxahlOzzZmaX0AFTPIaDTGfGQwte/fvWsvjxj/cQxISdHjgU681y1xj7HOBpxzIdJD40vB9N
wSdBce7MNMkVsuCzzdGtW6DLnrDLiW2MOSd+XuCxLRvXSiYhXRqUjUXQztbOAeuNhnHGOagXHLRD
2NuvRR8A6FgtJeirWYJoNKml0qm7rOkLdLMqD6spQInGRrG9Wq6tHsq8J0p/lJAHC3ojmis24gXt
N/0k79ozV2v02aIdgkyMamLmaPEKvBnv4Zpfwy/LaRvJzmJVg0RNM+M64qEqFTmhrO38BhH5Ihdr
S3S+XWVAIfwXEK+MNpTdFSnOCDlryJ96chW23ba9Th/TTc5pg5HxLvG4bWZ925bt4TXL61pBdG4F
ViYNxf+NI9k+MeSa2JDjvjGI3N6u3I5T1pn9eAxnhF9yk5ZFPAASEE3d04B8fUJ9ZUmj9zZTni6l
5zdqxeX/Zp8dnzRBc+EVAyzxSSoHN4cSfMNuIWJBekZFfUbTT9ZVF3XyPz1ASD/ZavMeeUHq3Xq7
wcSCJ0wnPTH2tygc25s3UZtqDK1QvSKk2mrINWpEvOWxilcA8iV4ejRD2IzrBu9SklhYFAa7c06+
ZBiz5uZC/UDIeHGk0UFt2+OqeE3c+u/r4sVJ02VuOji+HE7EsxLesjJC7W8NeL3SVURBXO6aDZ41
fzQkuiFGARnkNJC4XSnPIPfbzhEGrYeX1+FTwkCFZw5g2s/eaq3BfEadiAvMNFzdGrp1Qd4w3NCC
1kWFc+1LeraGrpwJheokm4ew7OnUX0Kx9HVVxdCi+fcyTZARFsQTUKl+uIII1snKqqM1IaHSoMBN
SEIzqdbvYkqLKzCWE9YY5pCP6MJsVFuNKCx7uj0FHW65ET53kp5av1x71IFvDD+u83GPuI6WelfD
Bl1UKcUS5LxzlAMgq+aEdew5JAH3Z5ewjUq+JLHNMnBp5sEX7TM7bDuWKN4qFZBQMEz6W3/0r690
GmUf+nkTjk0Pe6khXKgJrKkGgjfNcUnNSIqR1gRu4BYp4u+78vyCFsf0W795CxWZRaQTvN9pjMqu
3Bd101m1Qerwx035qAVELnA58UiriBCjaRQtywOI3SJIOe6xg6Zy+Ic0MOzgUEPdIXGpqSoIq7CW
YK15FjZVYdGlPJhU3182tjk5jxCZycOI6s8oOhkxZWgUf+c6luupWoqexzdrr5b6Sf/QYL/h/2CE
kn/jknKzUHvCLT4qBqYb9UlR3q0ypF8CPxEVxIFCgVSc+aVGHtg7rINHXqMaXL9Q6LuXPqqZooox
pLJwRMxdTO4NZtY+VufeYzlicIId/YexB+IwpgYcMTMA8LuEc7JGXwU8+QDBOfXcNSOwKhY3eFhx
l+C+ZkMZwBv0N0KddlZl8GXXdlezpFv6z9nz0CpMvtRqM1bgg7pwI3RCfe6CHYn2O7VMqIkeucUC
bDFNJlO7tTeNju3yc+Y69XnS32OMLp+6Tnv6NKtCmY5jGn9aWSjDoc2/f05/Q9gyDfmS2uTgsfhP
T3RpOR2zFNF7SnC8wmSJmHwZEEi27JppzWT4p2H2rZOtB0ZyWSYKm4D5HyB9CuwYbtVD8iYFwMMC
tpwFn5qBf54+AIEa/fFF3HWaC5bB4MTp+ZJg901Lcx7EgFSQjAmrNLScLkObuY7JV7Wtjr8SEyrP
KINE0N4i2M5AADeD5SgJgDCrDQHiCVXH/eInFGAoVSf2+dp/zNpYsc/BUsyjYlKPfQPhPVaFDfqZ
fjdgVkgjRp7Zfrp75i8hiGACvFqB2ABNoKZiYZxfhxhDBI81UvHdvYrWBpGFfg+jn5+ELUyGw0S3
YJqIZOruRFR5yQd79ckXELoOzs9E4V/lu7anAkY/yDlz3QZka6uY9kl6ZGV4jpVRP7oMNdb0mRvs
GeYNPsPN95but1OQzdze3x2WQ+wcNeVG7aqohw+6Lh0eDB7WX/jY/6Rx+QS2zrjrUrQm6d2BvEZM
j5YGs7cPnIZVDqgJ5PalVoV1sifQ7gDMCMxgaa/UrkvhjKvCR5Z97RUOX8GisE3ZKwGROatgBs4V
pp6rJG/NwlmRd8rXI90gip3uR8yLV1qNbpNfqzqp3P8pFxJFPt/tEHtGvY/Op8VxuUybqMyJAUr4
DsQe5xvMbbkq8Wz5mvRNqdE6IRf3aplqwC+xSnN3y9tO3vbdHkwgCOM+7Ju/Fxi6TxwYWN5X/eMc
INIyMlIj1rU3Tq6nNLlWD1Azie3n7D3AV6wrRrqzJw4SN52oYugxi3RlgAyEE6eC8t2qVHbSmCdH
hWvBfaXU+1ABX5mEUyN3xjf8iLC38sXTirt7ecREgvOJa00WLQ8bstupfYTAWhO3UsSk5kntmlhW
D1hvmksGNMExbqeXMS7A/VFqsa/yWzxQe9TNxca4ea6pBD0fSKLV6evq4xsYtXEp2+NTJyrTr7UL
vPaXyjvIw24CrN1ZW8z2rhorxhBKGwrG8BAfIonjS0fqFRohRNsy/n35TSssbAxX3hU7MRKFomgB
hTjCqpF+GuV/d5KOZBdlGpQDxaMC9jwJtg2wHYAN5Q7OTxPbCZouQ6ZgWi65zk1E0Pzht9TVp+U5
YMe2z3zQ6ioXQPJk0CxoUxgKSb2rJNY02v8lQRHe0D9nrfGR3i/cXf9maOEQwQgTWTaLDpYENVfK
PohuiOBNK0YyBoZD+Yu5qBXmLQ7TY+cQRf8avYpCxuzayas8m0C9wUcUczZ45by5vXPvCjcegPox
GnIjOCDlvIPVHu6956yxKATFYr2quoJwjXemjNlI5kYZ/xulnCoZWOQ4PuGaj5hWcAZtq+7oStYn
vWG6GWPHxW4fk6g1hOP38dokWE5ZEiOcV61Ee0GjliJxGJ3GvsLdZn0IQzpIGeH/s9LxwaxZVSUb
kYHQzVuOSHdSCGfsWl4LaoD4q69HrC7C1BU7o7gfXbdrHdMiA85bf+Zq1qi4Wa5ayOGv+pevhSmU
h0hzc3CWE+9saJntur9ZNOBlIomfNobDx+U3GIW4p6nx2sjF5zTpcoR0xRAg3CxcAN4ZU54PbRZv
HlsCsrQX3AFUpu0QejqB0IZdI2jaH+z0jJJrW3jksVfl6eLhPYeUaor5dDBMCrTISX9jJeyrJLy9
gfGC4ODkCzKc3FiGU9jBfOE5/cPpXn4ST//BlDjcFsd0b79UNUZlG+/YPGxndI/eWYM7NX2NJDhg
anTY9diqWobSBLxClul39fjiSJSfT9XvK8W8lFk5cB0cSwS2HHz2eeyjH2Gs4a2PBqnEldQfY8mP
R5tD+RXS/os+lvMi0AyX3xooIxVlemNtBtFApb7h1mHWcSwhr8hqtVuxtp7JGzvn5oJXBGqXaYe8
rYbPuRtu+vR2yUwHi70s6xuzLhMVYPgtL8skstFqoy3MwSkRACAERS92fPpdGEbBKKcpsW5fliYC
I/DamjBV++k0yszoDgwLVmqFODOkayKcX1uCS3TyJMcW4rXltzSIPLFPXGJzLL7Ll1l0sqPddcSt
iauNPhUw61uYvVEcWIPQgX1Ivsf7OJSoNJElA2aINSUh0fmFKYDkQUAMqanlGEIXSUXhIb8xXRxn
u3+BOchHBM+vx1wzXJsc/ZBvtPErmmEyG/RDHRU+jfYnEyQlaTjqVGbQBqPwwMwXCV1lpMlVHNMo
rl7As9PIgretVXvmKgQGA1zX2gGdCWHQB/w75a7VVqx0SStElZgxaJnhjsu1YJ18UCzkI0WxNn+7
lral3vAAprgVJwynRmoPk3E8NR80PXjXzQIIHi3xt65/Vwgbs5Ue6WidB+8aVqPcEZopRUmaXEJu
HTz35OHrsAvW86Sa2TDFfq/2swZ5IcMEuWbSOqc9bFw9452YLnEFS/uoE6fq3cMEw+JJqzfvO6Vy
SYtejlerdO9M+jT3KQOIVkwXhMFYVbSB5/Xx1HY8rOvistVG0yoC3pFMDbjrwTtH3FzHvAg+AqVj
yziD8fqfllBcBOyUxqkMNtkUVbNIcLN48L26nwBwf2lZpYVqejN9uWb9s+Y9UmbBamr9kksWPj9T
xIv9jbepjWQ6p8KeTxK8cxW24pW6AwtIYt+Q5bWAAWN6uBB7gxmnCb8Nb5hLaZS13gL8/w20TK/p
C9fAofoQU7UCOWqVe6Xgfan1g9diLnrrifDiKEUsM85VIUrgSiQj/bhtmre5DUQVACsB7cxX3g6v
mE4O59/7iRMRN/smJJBo177ZxsAYaJvtfCHplXeD2+o1KThzAp6r5btqcwuYRrq6TnzKtsQkZwxr
pZHTopEeS3vWZrbyzNwiUkzKJALEQS6zRgbcKFQhcDVQyPMYa7rYJLdroOPdgiLv7spdFH3KUBc1
rYWEnuECLjx7EjiCFczTaOHXdrtMpiPjr4qDKZJd8n6Vq28GE6dTjawL7br/yeJM9O3EFPmRdxG2
K7QqxyveWr519p1JFA7Rgo81DEv+0X2hF19wo4Ivz2xeKIh2VSZMQtBkssV0LCbIR6fYe3+z0EHD
CM/Rwvyt6nXGKMXHG04hsrAsOgiBqCD4/5u2GS0uCNLOwt++XLFEm4hSx8Kx6TH2k7EQ5SCsxtF6
gVHf1ckxFTp4gbmcGmDp8Ws6yTQiM2wHh8dhXlHEp7kr007dsIWFWNbxKWDwS3EtmTm3oXPaEKT+
O474LfrJIROjUAfdYoctnIL0BPBS2ri+pKHEbHUWQYNxk/E1B7wC93Fjbc3RQhgssBQ7MGFPcVTN
OILvs5CaR658HhPUE18/dyeA03QsG7fH98wj61OLCIkQECuwBlbo0pcCGWPvSBDNRIwMjsf9WLHq
iOPT2+YE29BUr7LIGFiKTAJmk8okhS7qggtd8pxQvPUAig8p1vU/cxge5GyCM+TkM4lPKuGeqH4o
LfjQQF0QQaSWgwb72DrQ3VvTCbeakT7HPcY961aCyhJVj4P7pab2D4fJC2zj+hLnNy29t4Qq/czn
zcfJ0L7jwuOYjW5eNhU7GDYNyVZ2Lo05O7EJr5UL2wY1b0AKEV03oGJhwH853MrbIaZY/VRvlEEv
wLpBQzUZrs1zaXknB+32EqQ0qWl0mUTrhFwe1XpCHG036ZXhCqekFQq1xKvhJjAWae1n6W3GuSSJ
HBjIwEc+5YCK0I7XpA0FmowyVH+bBXCI+b0U7H2VIy2/qaksTrurYfEvRXlxywhlWgYq77Pf7/zC
qoOpv7IvImzxb8MLE/CBR+izTk1m2AMkSUiw3uUoPqGVM03nTjVllTpPIZcMnLvKxNw9yQGluTSo
jHt4qir4CLB/zO4esVLF8SFr8C4oT+EG1LQpj5/OO8CGanwRAeRPiHz2z8yrncLYdeZWupwjSv5g
rm7NwV36U2kLnpADfLukJfCcWr80kqZBCytnGp5X38mt7LoRGkp3s4SYNflupPme2VFY4jZDq/IP
HohIBml8+XeDybgU/R27ZRK98yAAbvQ0aM0dM+Lcon/QIO8SONHGTYdJFerjuehakgYsAq7mdttD
Af8o7ovqNCoitlOXBWx1rT3FTu6i7uvHLva7ioASeTmLFBOxKz2G9qeCIyz2dQ4PsPwGYm3w1Tap
/BL2x24LQv5h/8QzoTBvc8jkdl2IExWl649sLmEby2GUmoaeot3grsurtsm6jG+Ue5sw8mn27Mkg
dV7jXFYiJjph7g4wuvBgHmsm17ZhkCve8bsd6HFmyb3UFIQ2PU+SVZohpjyoZlI/20y6AGns6LOq
p0BxFaXOUlpEmKqn/9IPFOFfYII+0cIaKxKdXyTUIKGjmdFQpnD6/yQXELrIkNUYYG2I/qJ5KJtr
iksJlI0fPRn1ftWkwW0ccAchoCUX+pVMmu/MfZIIsPanTs1n9weE+JyMcExvyH2oBSaT+x74+AMz
HolhorJMtDqkc2lbodNtqcSyCpetUDCevBGp/KQ1PgjUhLvpmMQjlrk0bcLEIeYKGBlMqF6wbbOB
7VLe60kG3dpjo+zJjodukLmKQE4F5AxJT7GDjElNYP+IOupyUcs5TSknYGzNI10tNEe/T1vBSVVH
bkm7SwVzzRVqpsw6mDGPtblR5OAFQ2lguR8sLiqcJuywl3v29ycyejvsBO/ILpc8R/BDrLMaDIf1
EHCEWYSK2Vu0cvbNBhqVlpQ6FPY8HXf84PuMekquWylJObi1caUFSHyjQRfCGMokoDMcd7PNJlh3
VcUgUqYKmYlVRDVVIC44rwZ5SKJeQbFFtts0muessO4anBPFWiSfSxyMoYBsbJc/xw/Avg/QoyxX
9CTypUMG6Y8Bf3f1HM16l8j1Pue3b6l6bFotAaHFynSnpo+sdnsksorX6qStpP5nSg+5jb8MamvH
hawo28PGfbgwC7YkADAKyPx5yUbpDizuEHYCfYTONc6J1HTaLr+UT1yoAc4Y8pRsoK6jovV4//9R
aEtAvSOujK+niz8usV1ZAP1IKI3O2nFV1XBwHgeBD2TfhcnuCspzwoVo2Aco9spTPBmh86D1W/iy
rkbWCIYn724NH5fb8QGkyZQqwKjAWn2dsXGkR0AEHft1F46eH66Ewhby//U6GsHqJ4icCWvGKGlr
40Epl012xFIRA1YAxoVruHdeFX+ozwIs6HguEXsRs6+K17nK2HTWWyCqyhL7Hm3IWnqgG4bMgKBT
EWu6I4Z2nMTDZCbVFgkw1pPGnPy0Wb8eXcKBN+CDH+bUu23xQ6mf5AKR7LpHqp347LF5OwGQqey7
SyfX0UdBZXMTZZhnwSuXaLnaoIlj80JriG2VNUJZDc8ypHVO0tH1l0KotmuSd5liWkkcr42vv4Sl
Rkx3X/iBzg5XlvVIlRtSomlWxuTq6s/nuwgkUumXS79OyHkmibHQKEQkSDYGDjYoxy/C1Jmdy7vt
6+mwluFEwCbzlnzr6Qleg/9CbYRSCYtBwuOaOwhQNibIH5s0NRGvmVQ/7KdjGrO8uIoEl/jKWsdU
i9NjbUpjh9Mp5BPBUUWlHynFWNWpBSaG3QNFRWD233s3ITEPKzYVbqQCyyYD+CxiBsDYai5ebSvu
2826jI675DjNQA08An9aLVzj1U7mEXNarmh1le/HY8+xCAj8fP+4g0JiiLfu86O2KUQz4QEAue7h
a49ATAQ9UlyfoWPdwVH8oG0fSCkTT0iSq1zmmnEMiLH2ubQUcHwNMzIv8lUNHXcpzgKlcCjNmtrD
QD9KRs9y2ZkaRE3zGmAN5wxHjq+QPPBmGhKfdr5p6+2bBY0GtZCFpObzbHSN4RQ7/PqS7pgHr5Qv
/CFpmgjKpjV2Lh++Fn0tEvbr+N8TCA8LvIyeUwvLh9Merdmt5ycDWPYqPqqfjpupk1ytnyBmmswK
CiV4q/imAClQoP5wyZcwewc8gOVuvesoI35gqMvo8qs0tVHqZNpCwGFuv1eEc86Qu/bZsrNpoBx2
CMS36P5Gr+bPRxZVELEIMxjWtPNRl7U2oKCIQkEVAO9qLWbyEhwDmC6v7iWDhszB3/ThVKQ02mVp
OsazGYfgO7qLvfB+jzSEek8EwYbNPJw/3ypd1ANQ5Tgee6tYn4WJ+dQl2iG3gWV8Bv1yJnRm4gE7
C0g5ngdrvCrhq9m9bQOpc9+odzq4gcCWQXgvmDVlShySog6TMuB1HiHdcW60DZZf5+5/2MkWa6LF
acYVXbRLpjs/gfu80F1kdsnbHx89VsRdsvTssukl/UYJQh9hl5ImuB/nCHJmEblB0Elm11Ylaxla
hSUQae1VWn32D7u/2MSg/TzyOinVOLawBLHDYUnMnWz0Ais8sWlC51cYpA2BqAwCp7MTXYFG131j
84mIbo0nMpxjokQUP6Bv0XwHvOcJjjkul4nHi7sojlvNW4YLE0JcIROyPoJCw/RHuqvsFMIEGXQZ
XOJnDiTCmxaGPyRWk2NmXdX938ruKaSw8HwHcCRWfLxcSJTaN+PvvnMv092j4Q+lruZrlkw7w0SR
yONm+3XpfXEbvTEBarAd1OBkvjUFxqndHVYuMBWtMHYDDU0H3/eLxPMxegZ1JxBvQ4HpC0DxEF8l
YpxoRHUbevuqFnRM5VzPV7ULbXpjS7V6RigbbP/o5sJkhbWzhVKnjzM6/ZnPZKlueBVAkXrwUirz
BMQz8Pw1S/8OrZ2E98ffgjh8dGiL9jFJnjiJWSkWBbYHsDgeUNfybSINskVveSAT9MVuTc6rCXm3
Th8s5NV35Th/VHca8TMtXOzfZWPBZoImRZ7EJMbKkS4Zo4Ll2WzeOm+TUfYmgBkg/oQLNM3CiUFY
fKaQ0mp9gKnZjNQlbs61i6KmGATVbHCmjL/piV4NFGckuBkUoSkxsuV8s0N2dbp+YIOMhefc3a6Q
wH5EDf3teUWG6+bGXqPZSDA7gg9AsOC2Up/3TqiI2QwpRnv1XLg7cAGrB7SzyRinWRKULd25za6m
YgZXC3ysDr66pC3yDh5kfft2+H4Q2simvmPdg4X2O4ionWSoMMtG+fcYjdPmngUiUQCUESxAxtjy
/QmIXKlzIipo7MnY/AgHmLkatwcGkdK/VJPiG9MyxBQYffdb6RyVO7hFm+LUS9lWukiGsDoF+WNi
gW5PMSK6OTdtEtK6PrUllE2atS5k/5U6s2n10omVypn7PNFmWSPOn4JpAkD2S9SFU3jMHc82YB8P
hzvK6knHKxtMh7mVQpIBb/38LtO9F1pMepo3dWqnvpIIgb5DP6lZj0SGjarzzzqu2JTvOK5Oraj+
/UvJReR+buxK7dmsoN5vtmef9DPM33kljKgPUFe8sqMtk3NvY5ShMYWiNNnu2GXMB7DYDTFSyUiQ
BMzz3shTs7qCZS7tTI2z45+nvFRYmoQB6OY1Ok/ipl8t4wEj9kVZS7v2zdjaOtxEms2Jp+jBGRpV
e/w4ya0uO7DoLj2GluLlL9r+hW89KOclN+ScM3iprdSpBdXdTL6S1lvM781LYTP3kXX183VBODvC
XO92KChQ6CwtVqEXfhHb3aXgP8fONFcFLR4UMd6NHZdJR328/wfx4rDZ6al1SrwLdOXtUj8kYSQM
M5TxJE0Ef+uKBKbgFIuIfUzDbxX79vA7qLtzWbM5xSMr8Pp8G6Terd0lCZPdzFVTubLJwelWpGeh
kH06uA468YJWFtQTKDSv8ofI+m+l18Ze48uIa7zVbYYA+11NAJ80vjBDWVtM92UvHrvMfVsF/Uol
ab7fJlrPBaw4pAAEf9JnXRqALuEqmvzYHc0eVJ/eXmThu64LGSss/7dFxWRLVguUg95xeWmNtq7W
zyrBJ1HOfxezFrvCXC18ZYpHuCg2v7gqmyt8BBl0+V+xjto4FOVmywLPa0smFIwFRTUmkzy3u3xl
UVtTrZInARChpjmYmXDDljMigDtg0o2sQFVPOF1NV7ifyd/KzLwxVJkLqVZbOJuBtZEMIOKlXhKk
JHAlJul0Kx/FVvYzqQ00elk4upLCLaoL4sbFDYJihF0cb9bNnNn6xgApIa/Mb4ZYCYSTSKl1L8SK
Foxz40Ag7SkxE/RupeBRPEMQPQGuRB1nN5Kr+FZ6n0efNY50H77a9pT9tNhwXky0gNoKq4IsO0r7
KzwI/5dkUq4Al/9lJgTz2ThSs7Msd9ywQI2GgT2bHJktUTmLKjY4FgSG2HQGUOjGs7wqHAlZpoUE
xBgsz53KCo9Qv32EywwmOS8kxjxEelF4ebW+J6ROTT51XO/7wLdmCx9Vjy58mkL0S3mSTZsgyK4u
xQUdteo4kCzi3wV3qwbolosTK2p+PRIie5Mypl5YxggGbOJ4otBi1NmnV6FlwhZU968apY5kfoR3
ywgM3bjUU9BnQxQ3jPoPWh5PQns0GrKEYTmQxFlens7PM3UfxW6Y8jn3WfzfkocJ4gox4unlwVK+
pCpHrv0uFB3lXIiEtjjOjIwNrbGIQ9YHs3qREqXvOFOfIHpM5o6ZIW1U2niISauLq29dPDsU/OnW
cxS8+IomQJ03QXERYEgYPU6Gt5XQGrr9xkVXaFXg3cFUdUHEgGvgSR+MOUncfZGW0mIit/LPcXjL
90HtvNQAeEXEXU6uM0m43HAL6S8QDA9oU3aIUncWhzJKFYmEmzmHP60lyWGEbjVIpf75fsx2lIsE
ff5Cm9g5l4d1IiDOfz42fcrIJRki6BLMLr5Pbm9/XNDDdqYD+Zi/YudQ1/Snxs/Bw6dFgAPHqCAW
YQf1n9NfsIF3+NQd9Ky7gKFj/goI6q3flFC028aTmEudPjIA+QDh0B3/qDGoiGja4sCoAoad03Z2
SDm3y1gvZSwTvQlfaWiILSpgYlgSCJ17yI1vWUG7RelHbg4QxwcKwZGx69nOtuvEaNevRGsSitbW
IHhjmyxDkxPf3RIIBOnyoXwcTOO02ln7CFasSXtNCIwAAfCytZSZ7axcKpmY6QeHxeOaWF8LzCJS
jSysfm8mE529h1JCSaUcettts6VY6UZlgC3E4GI0MOIvLjxRCxxac7YjZKSQxUYikf20hBjIPf/l
/me9vz67uQG3hsFRyS4O598g0jh3OBWiBKZ0/OzyYPJ0HzocneYvOAeteK/p7rKPJHdnmisjcljz
BeUq8drbxnQfTqVE/dKlt4q5rDVPgYh0Z2wVS5d+EBRyDcnCnCQ+Hn7xFRidyKtWPL6/0yu+yiaP
x5tDOKtyPZNzgD2uV+F9xCFWH37T785e07FEy3va1Snh1biGJFJCV8AYZE9bwCbe0SMSfC/WcL8E
8u4wKmcq0ZUdmjhbLyb+vSiIxJzbHZ3s/umQUa89I3fpj6MrTucvC/NJj75WYL9oIOjCjEmC/IKP
mNOEeOfbkQGgwojPMHgWFOIY0RznVUCs9z5n4fPFCjTBtVHs9wnrRSOBigAtWiNvgtazowb+2Yay
UsVqGhMiYuyaw/o5a4Xgv7f3Coq6SCmOqs8Ioc2tsKiqgQuEiWVMkKTxLcIiwegHlcVs++iqdTG4
F8q9pw+6ybY9b3IhGcPX9w5nHmGeCXz1jsq1NSZrSW7AfQcWB/XeRPp3GBFxgg7kF63UrTR4A+7x
UbwREXAn4v5zZH5GoMJTBB/R5Pt9ApyfMGgjckFJKTafq4gAW5GOnmMSd4d9NToMiJodCIDzknPL
sUmT660A8COCSTjl4ft1yW5ScrjA9B5SkRk9qCM3VHde7TOc13oRXg5s+FaE4hKCTH580Kl3ReyU
5a3hMCNAhr4hem0ufgqLYaNWr/9e+voIvSlzJf7rNk1vhceTTCSuR5QJ8Q2GpKEKjnV2oIjmIRnV
A1BQRWq2Uaq9xlAXbUbzN9v2NIJnnFBSSDErH9R2lpUFS4X8onUwcHOSdB6fFUQMKhHn5Q71LRXp
ghxSaHn0BiLD/08p4dOZEoRXqp0Tmib9aQ8WlhR4Ngly6mw8ivgV0QgIpC2vQWqaPM1ThN2niuRQ
CLorZPzqBlExwweTDoOufU74jOB3W/aS6AOVR4oYezdnK5V7akFdGJ0rnX9vnweSWsG2g4FNisP9
NjJQDuqWH0dRG7+lhpIEKkWac4n+NwfTeSSdbdIIFZ/yCXnP3ZJAemgnB2MnsxoO7M470IcOJ4R2
k5N/JcnRuAN8KIlURKNyfNY6kzAN2f9mg8CZsMPMNUcWHyQavLlwaG5bC2iY6Pv36pOisOj2lIUN
SZ3Q9bSqD8TGkll5pJFOXYpHvCMfKMBltVVZjLJumas8mJ960vSTJCZzNmWp1XA0h2e0znxLUZrX
H2GvBOXevKfU1rJe9uSqwjr26+sn6kX7xE35WMhKWZnFr2gKOpaX/38hVQ28HDfFqbmrBNcEcD8i
47nGEwt7kwrIMN+opH14rshVmGaQipRUP0goOnyBnYusr5VNFc9t9IpZ16GGcIHtIUuIh84HFVxq
MKLYSEl5ZNOGPm5tbAP/G2e3iXhEf8xTN3/O83XVU4tfWPh8lSH7IUYQvaU639SGQV3nUunMBTzN
FBju8UKSDlGs2u8E4B6VtcMiKy62tr4sVkVUgM3oBSTBSz60ViIfqnl4q4trH1b2oA5U8IgOU9b/
RCU9OH/j7BPCm4vB++SVHNzoBb9O0VsmBxkC96AzYnlpXIf3C28k/j6nCq53E/0p8d4A/34jNmxg
HvHUBS/1Fix5OwpoU/HlOH6h1ohXxVrUUFZVgyDjATs39W4OPbc4jb1kX+qZg+C/ZkmEg2HQcjit
oQkTpfX+bbFPwcAjkABFuNKbIiaygd7lREObUIvsGMYc8J0Gjprag8CPfyiI1+UVq/6ROeZ1kf7N
hVUZKhSE/NhO79mOLXDjKzazm1reDdcXfp5XJ8i5CPyiO/EZ+eBVO2WT/tIrwFxaOyyuJ2/1mZMY
tVl9S80N9CjT9bmMXrrAHknGaDKPXidECMB89f+q2iCtQP3bltgCSLPDwHFwYAMOi6nA5Oa3bN/Z
iEcQoF8DrWNrVjWejNlmbttv77yq/Rhvv2kH1x7B5/AONzZ1CzsZOc4yKrFU2mh9Kbb3nxb0UtzG
C5t/S77BWfuYz4ttAos9cAtLSKPRN5l4tY4F3ewUotLYtaBcXrWkjR82FHJ5bn2pdiAJcKSP1FaH
71ZsLeC6jADQ8AtcHkaGqEbvxtxCtgxCpZ2dpKhlSG4bVguOIM0jU6ephX0jYARsHK1PCsQrO83N
VWDmLWMsHwCoRtvjVZgK+UIERgdj3/2YZ/+zdC+7SnzuYNRK0fDgB1gbCp7mV/hna/nwh6UFaLiu
47o4WCofWAAVdHVtOLlPG95xTxKucEDyk3+oCwV0FUdiITvsx+0zvp7sp59DzdZebFm8wduDhVF6
iFwyEl8sbxl7VaXgi0cMquIZcSR+rpAmRgWXDxgmrGzI/kG9ZY4BiMEV7+iH7DEkCE6ZyMbwewCb
/5z3AOf9d9X5en7vfU9aEBZBsFQ+xtg7/vpcLEy3ImCuIkpknnXfZ9KpL7xsXHG9zw5PEcqGQJPt
3JEQaVKzDPU1kJto35qdS/Tkxlro+WzvaaEknmNo/ouOqd5SHW4IihlxIOwhhvFHh4CwfsF7XMWF
FA72IhsCZmgcUHg0XGaJtheJxtqvKWN+9HpThblVkx7bgaqvJw2gpw07oxHRIfQ0psWwaK+es3yr
xpz10TLDjUCkEYiaLOoOypaJ2KbNINmQ7NznbqiVVYpYSiAOFZ330cG2yCaT9SlWelO/UqRqnGMa
FJ7nK5jH7QGjFQMopHy1jhGXMA+/FEy1IhIFfpM/KGrF4/ot7YxcwfZacsEjs2d+0cbQnc0tFLwc
EbIHsQtaD5SPYvGGeBX5ncMNlbPWFaJYSErnKsGIE///aOepqz6NUchBLYa2dNBK+hBUtxJsDi9/
Lrmb4MHuFfEnzD9TKg+DsCm8iO9LX4KBnbx+e5j+psrErQGQvwg3kLnUhxKU9nZ891xGaQlpCpnQ
i2F22joDNGLkOo+YS0xDLapiSwohBPesbaY594cNhQmq5SrtwXa7b8lJkoYIYwML1TNisucw1N/K
kpOacNmJ11FDp7t0UI6NNurV7/HZsti4piTq6e8p34b3TXayrp9u90gwe/PVObcuTe3stAPH9g3+
O7sTo8lH0Fo4o/h/6OnSGj2pVpHX6FKD0mpgeBekcR+2lIl3rheg5kACs4lDRkXw5Qr+6dRPkDD8
jfBQcWTcjp0A9f5GdzQ5LZi5SgjdXsbGHQd4Dky4j709qwmjBOY6gCoQK02Lxq0Pu+W6jQhjNiOt
+0Sp2taoGLPS3LLsmzUU8NKlQk+D8DeAuV7MyoVJue4CxvvuMtCvrggmcXruhCzN0gvosO/PHr28
tA/xdSxXVR5yY8/C4DDkjGLNXiwLAPQydqyOx41tIBABAWxue9BAaQqOybRpuJtiFIloO+3p8CC4
18Ro6A06z7c/phjbZkeu4B3hsFr6SH7A+E5V8F/Utx2AE1ccX92uxITyC8GZPgW2BmigHtjnnfVj
uBP1M9QAmBm9r2LXdSs3oAoITnh5TeVglLjsTnhu6K342gC16BEHqBjJg6flBts2BBLjwZ4FNOyG
pcl3na8jyTrkM/5TdfrKu3cjTKpKJMfzgS8rPssTKHz3lRxSNVW/Dq+DZLIFVSAO+JL1XFlqVL7b
pzmn7CIc92FGCSpTo6tobhZfITjQg0rN8VVWaqpQAUERCyLnhFBOO+yHRNWiZU7cOdHKTtdFuWtb
DBIjAKC8CUcpzjG/gEGKidgFYpREIwmdbtLqdbdYIH/Oqe6nSNTNTNYqvQ0SvPWeMBsy8JuFNfLf
OoGolt1xel65bemgDkMpA+oXSwtzBWKnTiwm69355zpcgiAz6WchDRv6t6QVgEU6atuWCQrRtVZB
wcnKH/PMyBeqc7I78jj2u42n4AxBdC9+Rb4BqRMJxWvBE+Nl+BVNdNZYvwXtO1OXC+AUZ+RLkTHY
kJJwl3Pnovo1BfR27/vnpsskB+4xU0M8XzQSc6/cKSzHRDpvzAokg/bR7ThhKbyb1KwWJuP9ySGm
ceAOybSTj3GppUGpCxhpryIPGShm1+BEPxeJlxspyXsRxChLoHGi3PhbKZqZrCmTzj3czmZErekp
eV2B7fATwbd4NYHxn4xnuEL4CLEkn2zmEeWCfII9oVnz/81uRM62RhT70kATlBXtXe3wbXFSCgKH
ElOkJgJfbjFVCBbh329bTUszfqTr4kt3AaAHOEoAj/Qei21L5CKH93lX67kTSe4NrI64NYn6Yj+S
T9Bvx/OU/zzZZ+lSY7cjfY86LAkwrEn0y6PW2GbbeLoY95fSSNUrgp3l2lmmncrowDK0fy2rQB0e
xhB7SNSCU9nkqT6Qzdu15eBVwMxp5F6DC+zfdMuX9bgwbAWHY0eJodlFGeRY6ZFatduRuqOsMa2e
5eZDVqaueWZUIy78kfoH3FrvXnHBTWffys479Tkw7N9ECuk9aflRVpUE6AURYKu3AzDDdFO6W2XM
7rSMOOFF5ytaonSK4WyZVpS5dMWWGF5ARF/YcefT0SodJLXhrGLYhkEewViOpdDYQuJnVUrPi0f8
2Wrqh24dStB8Hh4GRlTsj8m4HZv1sciY7Tw+f+LWgnVgFoQeE1pu0BwGXU5HJPEMlLjwRXfdWxjs
DTxfuagrmbAhQxCzT4qC2Mk722wxDN6Mk5vs6s5+k5kxvfRqbCEb2qP8/TP/YUGHWvrtIbFNd92w
3x56S0AVhgsWQR9yYkh21yCnqNGwplp2ZvuGyVRlwVPCsxouZQwYDuDJY2d01GPlEvlyvET3PzUX
O6FCRquy/kGaBg8LOyrNEfnKckmWqeGG0hdyzsVpTi1kJxPc+HRY3kJ0PXxlAHwHzEO1dDbVmQXN
zrVqTPSOIjcZ1SCCDd5j1pVy588s27IeO3EJ7SxeyJEdaQqb4bDR0jASZCI6GCsKUQ9uFYN3x4bJ
8696nUA0IJvNmPFyIaIv4fylQXaNfWADsS5wa1z7SENtHkc9Mm7ijNfbYmZWdXUlfKtG9aZeeL24
ORMuvbWA2fEQBXZLWFJo1OHYMTDp3x6GC80JqYE1gLH9Wv1UdjrR3WHT+UnkB1GPhn51+OKxECgy
nTnT//5tSSjK1mQeyQPqHumgxlAU3GBbMeK2A56TEgk1fJyn2NAnV6fRDYw6lZMA+eKmT6rOXpoH
Nz14MEGcw9OODh7fOCbnxQnm4HubwoVsdutRbitYTtXukKsyaGQ6mUMKU18Kr2yfZuMVeJSfMxH+
3n83yM0AdGcBmjvfr+xv4bwc0ZDlOXed0VcJY2gQ92kgeq0qnWzENF2dJi0cyPgmwqjmx0PXvzSo
C9BMNnaMU/ASCV/mjeWAOFTsbsQsO2VLmwYrTGv24WwsirR+AfnCC5HMWtTxT7JML5H12Vva0VrX
tJvO07iXyEv4cer8n9cUSLidm+r4yRFGaQoRYhyIxe+TOWrFmkva4t1Pra6bYYTFm4jVm6ZzzQIq
3QUpQAzHieLSs/r01DX7OcFMV48X0bGjPqPNzP2WAa6gh+uCAQGk3HfkTE5LgLt7cx0ViXuYMHXi
x6Qw7IHOuJ4GgAGEmNxQQZNu1QGWRmu2H/y8OdIKQOhPI7hb6c1jNS/DZdjc5jVX3lzlklNPlxyy
AI6Elbr1xhxaWh/wlxdgwHuUnV3In4LAaGUMHTcXZ5RasCyzG81qQS05s/0vutiks5omgXtXNJBu
cNYim0InW6bqyQtscQ5CKWeAcOy0w/LHiaqyM/M+Om1vLjO94Yob4yTtEn90dlEGXv7AEJKbiUV5
O8ReZ5Hv7ygB0mnMYEi5IPpOo9JoUtQEE9A4uPDcj4TPOnEiM0cmspSDori1icCTr+gi/W2qbfti
6cJUtDmdzz68Dsl0DeOuqvqbKqwBIKkH1oJaCH/PewJuCHqkASpieNDBMLGHxeQ1uPwX++earsFk
p/AP+NjZ6m5X2430Piy488y7DEc1Tf7jvWbvLMX7gOYwG2au9L/9Oh2Hs94LSWRaLOcaXaMGF8mb
o+W05GO/fTzZeuL/nGHMMnMy4Z6hI9oKzkjHgybhm2hORdUcwZDnQDAu9C8OiZOGXpqS7E8kH3mG
w5PR9ijT3O5BwiHWucfrTwxZh08qEspeoJG2oaHnzEZHkaG0hHToE22X6BCApwAgoFAZL13d14x1
F/HgjhYqdH+pSu3n6de/fI385TKVN2nH7zIkaxHrwBTjKyyQoE4ZZwvlkXWzfZN15cEukkav3VKe
TEZ6HFRYTmTiMT7zPM3L6RyapWoP8nQt2nDcXz9sywkMW1yTPPcjVGI4Tpj2ZJbiEqoEaDXkuho9
3T4qyVF+mk0VTJ4StGaOmtpKdbVXX10Xb5MQOY/5MwDoGh5e/tkMdu5x+cn13x8kiCOAi+6QHGxg
NI9HlIPA5ybWKTDt1wSwFV7iKr1/N2Cy12MecCaJR6PyrkYY35NsOtQNNPE0vqMkhTH/nNhpKg7Q
ATnuE/bXu3/oNxFJODnPkKVPGZzsuR6E1j8qVGelfD0m5X3ZXcW8jZ6TCDg9+81Ha5ZDJvVwSkup
b8pjapjQBdoHq62gtG42MFGDS81b0IY/pvoJH8nXDPfhUS/bCvvjjB4962UleX5Zs9+YH8C51TeG
yX6yiYRlhJAk9qGgTPvVYak2FOQb+DT8CCyJYV9i0mWn7FhB6GOY1A+wV3czt2QyiS786EQeS1dE
jdZ3ALUnxvbjYtbnP4YJCztzpQrIenA+shCoEGGKqFo3ZoGkuMaV3wg6PSdQYq/C18yZzj29Xi0T
outgWszKGx8ilX+bWTSerpVOVJwD9XDyLkz4Vt4rPWkmyIyocBqEVldKyyUmNMak9iJ2ROHBuZf5
WwaJWMKGp6I+myWjyDSqJk3ZW/i5l/uL0C7AHNlCY5a0jXrXMm4FgDbTE4f6a8CqDQOd1gMs9CNC
vgBlJgzpAiAjYKt169/OYJx3iKXfrLpcuavf2fgVN26cBraVpAX70sKrJ+/ELmJdbcbhywyV/gOJ
yeKNG5ZPD/bF1bAikFLkP8t9omU1ksD/y/u5mzrUEmUcD+ZiRQRBRZXikJH3Bfla0KJNu+TSwFKS
VAS/UeR4JfHTDxPPwlR6Ag4Rl7vYFvCxUW4TUU04+lClxx2s6KV5MFJGuUE5K0SgqIvzYmCT5nCt
Lu0hH2z2ZSfyGEj/r72KYS7Irm3/hzOizDafhqnRmLKyamw+r8TTJbaXubBEP7bmAPKrjidq1GGb
oumwnNoPiyQx4HLWClIcWd/tItw7h9AGy+tzd6S3yG4HNxdzx7w6IZ+yp8uHpKYyHiXw89V1lvBy
/Hajz/HxwJaFgBmipQpCVf5EeypUrIf4QwXMYv7b8+GxNzbBqg9zRHecdfFZK1wlddklURiWX1aL
HrXT7X1MJqrQgv/b9NTZ43LKxs86ULrV3oO2uYQrcr1P7JUuto1a5s/d6ljGNu3m81uu36YBv3Gr
4behNW8eB9PfyFl3ayTpQy6Ru8iz2oE01KLyx5TE2X9yVB05bzBh4GpmmEI1goy6tymM6CvSIQEg
hjGgFKQrFZqFKJ90AAiAIRnW5zyjlwzUTYt1FUj5Z8xbDVfas+Nbc4l4GKtGTy4pf//9BW21/YhX
Mtl3BrNgXuk7KMYxculWRfjoB/b0QFRjc2mett14YzTVY/6+yT1uk75PM2OzBG6vximh/YYviqY8
jSGr8SUx0VM1UFFMm0g5C57DBMHm7T/KWfFGapH6NOzQ9n1kx9xRQs0k6cpsaoe3ANA/NAKzj+Y3
XO88+j/9I8UsUiZ3ngNH5GugBFZNIheEYfs0J3KO3geHrr6cyO9XS1Ca+IXr0lRTBN2nxOPkrMi6
xBcr4BDzGDub9fr1IS3+HLu5zcaIfamu78CHch0ZxfSZoGG0lIVmhjx64e66/fPQYn0cM6+cok5W
wEdpzuK2F3Hrvlptojzb49AFAzvHmJ/LAGcssdCX03ZhHUL13ZSRpQuVgvyCDMpPml1CpeBXIPZS
ADj5rOLCQDlMKyKa9dUhRp4O7Jk9Ya11cS7QeiBazHfGNRx5Ul9IfBqEwzo+dMWAJyNDJZ2fCt0E
sGfDBEzSQnPhJBPAwquG4awWoCLgfPgl+8HaS/+Cb1NdBdfmMRVJGyB6ookQ3mxO0zHbW1sYUTtF
Yz4eJYtfnS/Rh+X5ySxxOjLc6b4EMyCfXmVj3/oPb2j6oKvbP+hO6DtUKlz8AepALAIO6Mu709Fs
jc4/SPr+SQgW2SMDcoKuuLbuVqRJKpvvHvWyEwSRMEDwprex2F+MaIMmdxP2bBqwshP5W2FEldnt
Y8thiKBSQMeo6+IrJd9MNQI85ojb2UchKVBrcMxoz3H1r7cr18ys9X7zCO0I4aa+j477jtTy/SY3
A8d5CBeXWwVE3afbAX8Cd67oSSsTu0ifZm32uc0NVPIh74SCRMv28aRiLPifH/CSbJ865H2remvq
8Q6pZrOpyWIEUnrU1HjRzqjBpYhMYN0XdW56Cm6fy33E0Nz45tIQzKpjUL8vXoIf4NjJ61b73VDY
zRrnHCeAVYqHD8Y8bVsu23812fgj9FJqMy/P/lkBAr/ENnfnDfPFAT0SOZV71sBLnrGzwUxfY7q/
i+5ZUEh5QCpwwKGAI5ajT5Qkui1b+sigoXZ90uw1k+Zy9UQGkc2UQz9EJPTcVed3BNe0Ps6qWoti
2f7DCsSVsyGRDh6KjQM5L9yMSVdK1PtPaorBRSntqK2Qm9884TD2H0ZuV50H64kOFZ+1utfM/gu2
AQzRHuYjVddPfnfMC7y9Ku6TocE8+/0JqONI2O/uh4timZTQbGjKSSxt2YtJxmLpPJmycwKwQcBq
7wN4uFVXbsTxoBk0CMeoRRXL1lIBMlxkOJshqURX6rUbkVtG4lhn2i4c/Ru9vHMuxRIxd1u7JlYR
KUXgZ1i1Yx/njmoCSXhEpvONNRuyE5gDhodwLtVEnyy7I4nkoi5uRMbIo1JK7CdRf7188r2JY/+8
Po3HKMHRfiZonYxk8kxa9WOscm6eAAN5wTTawpJMTOOiQBynlYfrUEI0/Unpf8+qhNfHjCIKUaGm
BcJJWufY5EpY3rcDN+PybDE3v86rFlXqfsM93IfZQwsj8wDri1dpDpC/1wTwQGVwxBuDZXy5FBls
QvFTeNtxUTuxDThYi7pCHFtNyMzGPrbDzXxCH0lcOtjy9DH4Aiyjewe0XCyFkgVbWgMBWASasU+o
GiAouu4mCJ97Xe4z9PI2wXHlQnP/Zb/knj/wT0MoxEG6ueIi7HWinqZ2H7NY1pkp+TzT9B80kFgm
7Dh6CPXOs7Mkz+gKQ+jafO+Wkdqh9FJHMMYz/8RstNSIY4Ujgx3Ge5heBh20eUEllICkHXS5P4tt
bbVr5GmLW1emdmvqu6M4+4UVaeuE52vMWPo/zokCnp7F8aG0zm6ET6bGpm2I6trHUu1kRWVXCb4B
9YbBp0BM6yLh/pLaeo9tnr/l08wq8L1cJTevxPOaN/5EuyncqjJ6RKZ6D66bP48XTYIsXFBYBJrl
rOkB7ZFfPsrSktUN6UiDGaAqy3Tn8SfBBG0NJLpgLzAfg7GLwf4ruFPhsH6Kb7xkjS0MIW4ajC4e
ehqkNQL4xzGovHX8REbQ0fBwsNG1TY2Srmxov6982NodzfHVYyGfotzSXvoXAIEkZgo8sDnQDh/k
QBiBOT7QH4CbW+oiHzcvAy45dsMK+EY8FHFD5v28q2Uk9Qcg+eCLHWl57RQQq43MBhdQUkJIYe32
ZIm4OktuI9d3PF4KfGH5LYuIIS2CVhaxJv/688Uopq0kXfsTHgmGgSBUUfmbsmEFvc8joN7ztqF3
yk2Kwj5Q5+P5s2ukdQoiht4eTiEF86EJk1xHBxxxYB3JRekcTkwk49Cujxo42+10KlZ4ntYrZl62
6O3aAaCS3mZUodlUIqCzx4VOctnFubPNo0J4N4UYDJ4h7rfbN07HSl765kyjiy57neheDnfzbDJU
gOcQIPF0tUTCN7OgkpAOxpiQeZiDizjdZTZ1WygI/wO4WonN8GQPFYzLiigmkBGrAKSswtHA5cRp
ZEjh+hmiKMC6/8N6b7+QUnMOq/CaFUI8VQIYxMuN8AZajrm+SyGlqSXmBgqLEsYIPE8MXgZUQ9AJ
8XKKyJuS1udxEvZFj596r1Z/R6IvWpGP7IDlKi3sc7M2eBDdLi6WHrJchg+ZOQV+whEmrf09aV5o
YVpLvx3geh8ClovzNssr0smdeGI/3hm0oxsKTmvQAMUnuDL8gUaOuwOEVc0OH0kqNjKpVK7T9Df6
qWsam8417XnvIrkrU6L5HY84fEDEvg8TiIRnigOcDfTW+F6/59GyWyyKgmG+RFMC1zP7arYA+dzU
Nj+Y55Ri1ojpSjqeP0UTcMyWOlj6o0ff8yxOq+7CaQ9JTldPUjvy4FU5O/bR1eHNhMk8hpF/aDz1
MOccWNSmjZ3Xdy1Nj4mR4GD5fWZsiGvQtmY057cGaAUQNFM3w+XMi8jG3p/IMyiUJEKIjlx8qprZ
4NuuFzWDQb78yajj7+bohCedlRLWvIgI34WerySqVk6yVjUyow/D1cTMtcOoTNUzsDqCp8XlhWwI
3xyhtc2rspHW+hGDT4bGpEZ4VVyK4bza1gejtPZDR70eg1ti4EMqwdGd2AtFIqxwkCCK45SEwO2m
dJzgF/O2EuAGRB8WyfGazDh2JFqbuk1hP0MH4JU5F3iit6dlTdNdELNISXZtArTKxF3KLpfFWYEW
amv/2ZeLT/GMn91W/GmM+Svu2C74os1XL0u/SGk4MWvVNZ93YU1fdthcjR45G6Um4PQblltOu6Ac
AzOBnv9aXN2g6zcNIIT7PC/DDRLu7h7tT+WkQ/+pbymmL3kboBC/+7ZiowIsfUWpSkYfmD0rb46V
KW/DhO2wSzoquCx/ES9X4G5HJkW1WdHWhfTtoA+Hn8NO1CNKnXQDleOkDCDJEamLryGhVl7msmL0
3y6bjzZSQMb+zhR+T1ZET/kvdDoTKUipskE2p+GU+MVpphFVqBwp/1NAuKzFseAi3+afbV4GEvRr
Mmw+EBt90T9QSG70Yum0fMb2v7cCwKcWstkchP3g4T6qFOAT8Q+HJXqklCltbEatTEHqi21mIsav
XrxbxwZgdpQ+yPhGd5HCGTdfBHrvXLNEI0uyRWQ/ryK0QIDBVqYyDUouUD6IBaV/FxARs5ZZ64B6
e9hHjnAwdbcqDPZL2lCXOaSgQeekZx99TcTZPYT2b6xkxibDbPd6UKmDMqbhL9N7+7yOu440ce6E
IaCUm76c/uPcyubxCIIAZqfJlWHZO2gTealVuUupdCM+zOE53Aip5Kr8baZrZviPft/bzU++7Zd8
XWBC/kdRTy783bpScWUQ0yQdJfK49s8H0q5bYlEGQlLHAQj1wauW8E9kGpwLMNug6TlFJmksUEVh
XkEKt3ZCRSF4UgdveGzxE2rGZXR9b5Vl6h3CnIoXg42KQHzUujqT7Z/7R5cP5ShPN/FYTXOv3s2u
OBnvnKijGWgegjor+eZGcOHPvZY05amBGiB6GGEddPPdboUJEF8z6Vgf1SgiSER64vZYmUeKSay8
+BrPG8dK3TmMUX12LGNc/UOFd5IQCHa7NcvUy8xTIbPGxQqRDaAEb42UWMaoUpdV1BYbouoLSUH3
6Xu4cXAL/y5IElQocF4Q8S57ZrnwjOKeDQT29YgLt8/o0/8BoboKkt7Iu9BSzaAUQCb0nO4Ikwn7
vhoJHJi3O+eXNFMdssz3KyNykB4cupKLOAgoQFYIslJKh9OyHsn7EUzQabVGY2+tzSRxo+ludLTB
DOF+1JJOLqBDlD17R8xFRDByskAyUte/NcKttOXNexzJxHmW+0vEkCbJU9vCzvCqZV1b4KgkpsHI
tLHK6TfLxGJJ5YDZ28Egui/ZoByVRXySiTX3LD5x4g3tbRr77FllLJzvu2X6lwzmJTRPer90oTsL
QlQ8QFFAIz+aQIjzGeojI9k30Mbinhk7CQW3zaDlAyASeEUp+U05FCSWr6ba5P8Eb8hKNOAEDzZU
Mp2xw1ZRGX1D4ixtExCyFHn/ST2f+3ga0fILas+pVRWJi8okRJj7eMOozV6y0Fpxsdf+4kG49CsN
f0louthijtrH4SOBAFPKsq1gdTRz4iW5LNSx5hkA8t5yylsaxWSh1di6CD+pmVlrsWefr6RkIoJs
iOSvQ+kBUoRjdw/yCcGmj8dPI6jlouhl60XbHP9qOd1pOdxABqgoA4fPGAe6MRCZ7EFd1a/RNXGJ
p01q8GxFHvaxaL7XkjuTTFpcpzDffWs+Z4MBSCtE7LEgJAkGmyfjJnFuaZAr3Aigp5dnr2a4bMQX
7UucSW6xEUvMbfQrgoR6LpRYpfu/oJC9648Muax7mjcZqmzgCIgRbTe+GAqyE1vGin+x3r7WBrjS
ZDKe/z6SZSA03Zy3bFsDBzgLKkhsQQqnEg8vKmBiDZJjd5TubsOvGPFce2PslUCPXTyVOs5IhhXE
nbPqaX3NlHF2iC+XleUCOVPAIfoecfFtCEcH4brTW9b2Ncqtt9sX6EJ2y2dWxTLvWg/YWAKEF+Fg
R1aO9u9Icd+CO5jzMW7PsGtW07CsXjRixp/eQYzbKYtf8Xzky6PuYDuCCdMQMhL6F56rsU71eHKN
BZ5VU30Um5fhYSweuzWhGWgugLVn4xH5eqar5ItlbvBWaT6nJ4v9b1o8dsUdzfLY5XS57+tOqD0p
LNbKlv32uzsQDaWPJVfHknPSm3Kyp9g/1yQfk93CIyvbdUjO3ngYM8RSH+9fdKO7hc/3mgkN8vBo
79hwNEb8oKe/rs/01L8TFmtA1ccsVIzmLvTCFyyOiN7Ihhi8Sx8mORMSueyheRjvIB7JQhdRELkV
o7LY43JgdOuKnuWqq4gcJzYyWPisShcmZeMcNSBADUOvlfMpS/xA7Ph+XxWv8sKpIemEhD4I+iJF
fPetW4+NTyVDB6InwjgE4dpENa0spQMgD265yRiI4HiHt/YQ4b/Xf9gBKruT2g+J2NOkaLlLB55R
KLmIWPMb9z8C5IfP4kqQHSPzJ2wMKkFhmCEog8AagJ9zmqEhZGmctMdJvAEoQY32uxbEsooAX5xF
7IpyXwqtNC5ED74L+Q/9STi8xcOhIq5ALmFbX7+fPYAbw+OxPMsgP3fknYuNgPR3lq+cVk3CHK/a
yrXXZm2VoT2ZIQ04p20uxpgksxuT6b35b4bXOKurMluSjk6sDs8eXPg9DCRf/+RM62+eHCA3FKJ1
Da79iKQzolxj7zLk76uNY79YL5vDVw+ItKVnRcmZTxU43ZunjUmvYwSx77q4xpTScOTXKxVlgz6e
Kzk/4Y0fXMXZIFN24VO+ZvHRzKlwG24CRRUPv5WPIRXgcC64Vn9FzSOXXfjKGMxBgpOMK3Kw6p1Z
/eUc0lHcK4/bbk/5ThUJvOlGvnNZBh4Bd5OLjC80m5aoVUrzI8sxS3CXYovoyWa8I+tFfLQgYWHV
ccojEBD4wlqYzxAJMPc7quPhZkYyJshhsXWP/SVIqaE250Fx6diaac1Ta7NpJ3PraJJM6gsnPXpA
U/AHa19A3l/v+tbQF4gwttDSRbNjfIXJeOorn0PJEX+c2OH6PW3lw2Ycj3kcTCkX4TAskr7B9vMZ
gRNEs8Lypv5DSGir4ueaEpgPUhAMva3x/p1uuX4uJMtavtqaqBHWwKOrObT4PpKx+u7ZGeM+jszD
uFPZtWU4sI2frv0Ojb3LNn+cFL7jkVYwxOU9f2BzJrI0DvsjUXNk+EnwgjTQHvMiwsffoavcZDOt
atM6VLKra5goWkHDL9C35y4+M8Jd4zRxsEzLaF6b9tm8z3pAY7NL2Bcp1e1aM1LTvVNa8nyE3s++
RDvEXkpQ4EvCBbVuGJKzLbvQISAxgq4PJmXAQRKneSEFloAu7j/ZOQ4amzKsTcg6d+Q2oqSjl9Mz
DJpex4qsbho5FzsWx0cGCgATzOYvvFmPXL4gniN2RO2hCmuWEXkskAtji5A17B0YIpBDYwHcsWdM
v906OOiYoRWcx7XOwTt9T3AMo2kEhlHHjSsHVi1fWuoVw6hH6UyZbmnQzkpx36TDaM5IAwqT2PAB
zKa/+eo94ClD7HMA+wat4hx2VEe2gAXdikREM+8WuipWzjsHSTJb9jcBoZY7GB5oJvsdB74FFz1o
+0A7kR0tKznTG1QoMtUs6Cci5KXOW3R+toCKYFs1myY6AyWV987k726IM97aWnlkF6cVYrab7yRc
+0y1IWm3CKACSQVrXxXNg/fVFbWUqbp+OvATXT0YET9E4T1xZnlJrYzFqjDW2vnrJoMQZA9+h4iR
x96TX40DN0pdLuM/1eJuFVhFE5nwhqJvbd/4BilpOrSubC9NhW08vSm0Ue6t/HfyoeMRX0e6qfmi
gmxbYbKc/+OmiEj2zAPAj2jKxjVIm7T9hvdyZRJxOOPv/G3j8sQACJgX4+IMFtMU0FV/2/7bU5mf
isvlwQTphcaJV0BP/SH1SfUqwnbX2KzNeVILlhL21oMTGJ3ETNY9GPFgM5f+HGHwCFf6uJFwAXzU
HUfqQtpLRmzZN9GgRKNOMCBJyd8bOhi7KYgpnG++a5J4nMlZWb+n84ub75k6/jdtNXKIbqBO0NsY
q6+2C/HxyYNJTLi79H7qA/AtOiDIA8slalW9GtfRkDgjQJafk5NiCMHf6lpu8enLzsmmLV6RpowF
+eZ8R8YvB+Zu3uzxm+U5wTJQDhoypLFdXRKpFNMVeGlZnM73GDknfkKcM44fp1yX2nB+KjEBLp05
DFlEmVI34RZrcGUhAJjZFMe4xAN8PHwB2cBbZ0ZzKVycYfXP/SCmcCxiYTQPIDzwhIMys4Dcguve
h2IiA/T3YKzKttiSUVdYIVOGoEM/LvzWCyiKvb6NbssIyoL1x758IQfPBmjxULR6VV+YWA8cLs3E
TtiJA4U34f8sOz9OGWUbzmS0NGDGyV5XT94QO5u9vLRuqdCnuV5+Pl5a0F0w3jZvqmeA1NB+h6j9
gzm1FpVvrMD9o6pyLxdPhHNFM/O14BoZ9oKdOYzBuF3J9rWZK2BHgYzDXWbwohs6GKAmN4grJpUj
NMzdlKveVHWpMMuqhDEUap5cONgoi6Vvs9wX2DTvwhwwMptNiEoO8XhSvO6AFGTsYRgEaXVcIPRX
sCbOqQhSqQJzf/c4lQUY+6zaB+0ygC8iNbCcWb54bebWGqqcE0y1AIcfKdeMr8UpdxuwOZvZ3L6Y
8iVeDA9T8962s2ChJYrj9FwrlKT9oJdOOqaRukq9O9+3UA549ptWEh4V359W98gEH5kMbGn2gpTo
9ei9nxJEt+r5geotY4IFfQui64NDFrb9DGLMfDJXP2tTyfP/WURk+TmjEj9VubbhgCPi2spS2PcP
h+CUeVUgLxM1GBHUoQ/PfdjXCKLbe5Gd43UGDdFq3SNneIV0WLnVDyUjujdjsdWE7bARs9PNXoWx
DG+s84+Whk6aT4xOPUAbdyhfqTsJmBAQQ76W46qfpAkTQFH9OSw3gAUZMkbg56f2R3ZIBXh8imQV
XL/HwO4aSCfpW3iuvgwbSZ8Zuq/FfLBrDUGHlFTWJDiLTx+Sp8bwon9AjMAN6eY3wPWZGx1lQJA2
PjwNiqw2lpIXpp+zbLA5D2DB4Uws8PUrOIHN6ghlxowtPf/0DiLcqsMEjVS2ToHFiM1FpVVVmcwm
lR5CWxIQPE3oGLr1/JmKigj6BMqeI8kkaxrPWu0dshnola4T6ZnWLrmuevs7mfHXh30Xf9IUgupF
R1qq1yp31tyG+CinJIrykB7vAX3tvMcGCA1PSpLjSDczADLNpkvTlJ6GRG8b/C+O1YOdKZsPafdq
zeMENYTTu0iz3+P/4RlBcogwU5IghBSJzY9V/8y9jpl6OCaloHnnblC4lSqojE7++OGFKu1G2LRW
5P2DqbqIZtMU20CcFm0n4cEnfrmJSlaCSw+KNjKn3YtdW8p0I4q8kBj4g3XKLdvmVeQnwXrbFRfy
BqcDDXCUB2VDfFP1kt9oRHwDAd9H0V3ywC8ZA0FGvGZcqusNM8aWKhT0OTSi6oBDESQ2JqwKy09T
/F6joqRRKxmRle+vda2U7KbyrTBMl4Er0fyf3iv9wttVyaQe3/qN4AH2AWgL+Wg4y0qvzG5Gf9OX
H3ySuzbUB793kJH5TAqueYRX6NhsnbfPPx8Q3wJkn+MHpZnzCLRrfNkdclwkgDJZ3rqMAeoh/otw
TUtQOkLIPL+FFWOufVAiaZ3uD+to3Vr5kqzavdW+9aeYL0XWn5C4mEXXAXTfYzOeik/SNHeXzMf9
ZTFpMK2pcBu7tzy014i2dBzykSwTsyPFC/UBx5TeKghz7q4RqRxw2NSRF1zeWMD5B6s0d5BD8b48
iNZZkJs04AeaXnQW57y26+Y/iUDK1MGvhqfL8OXox4Gi7y4gZqT5bVqkWCabXqB55kf7fVXukwUb
f5Fh5Tjo7JjXTZWbiKsM7FoTh7Pn091W9wFxBjJrUhSO7mYgQ3aahuwlxqlFCdBmgglfuSxiPcgy
lW8lMExVs0Zk6n3JWFZdXGxyqqyZXxJVykhmBJbLAZx7leGyYQOCVfixcrlx5QYjNTiCJ6uViZUH
XWqNGWCENzeO+GGfmhkKuHmn3wIHH5RGukeUls7XshmpW1s2bKkjypkGPNC/+GRsNg9PClAeghWr
4Owh8Ay1y8NzHifd8Va+cnpZOSKh0Nj2YRukU8+K4NRUK6pVKkqfsdxrdgWCTSirBqtpx0arYYgL
0OvwzG7ieKgHnV+oN6JAcRkBo54P5ddrECJ1IoEcdzgY7hxznNfbE/8hKSLPcAwBqGU00a09DFQA
o4QFsxhASIYltmb7UmFm3mHim9pZyjjH+ezp89brKFIDnbKOP3z+N0pOPTZUMZS1ZjkBwq7hAj4t
VEpDrgPbtZwsQLJ+Ce+sO/Lvi29wwJeHGq64x87MAUamMSeeMivCAASoIUUoRNDZTGsDnY6bfayi
0gz+hUEb/roDaQ5jOOjTnVCXX6lJUTQ8v9/UUcXZllyZIQyZXWjgkWmxA6JGBEHP/KKvXVYIxnOL
M6sKD7yVgmWoVgfc4s+1n7eCF6ICxWwvDEX3VMg2VzW+S+lDc2GFETgRwXXb5lR18LZoOHjeSO2R
wIiYmKqvxn2cNp95yxpYlGdFnRnJbgHOH0tfnEcZht0x5CryV1+h57u1t2UyKgb4HrSAD08DPQ0M
q5WH2rrl62gxiYa3Ybg1ik1AE/NUfqh5hEWOYp2doIJZl4wi6DOTt+3IzOy9miRzrfUQHBMMo+1j
3fW1+iEUszNmZNGrYbGaeCZ78sXp8RONUEeKekiiwU8BbvG4n4tQ/pvkNS7sxSiAlPx1OT7HBI7g
RTh3pOrnrsxbTNOQIH87BcOJXYQ4ZPLbsiSgYfHYFP5uSNfNCVnW/2Zyo6+nLufI6nnYPrTQbE4r
TytXhA4jJzr7KpoR+d4Pi84g5K67EMC33D+K9WqD/EWjBghc279uUCJeM/reApFu1r+a4qK96gNs
iQeQyU7pYebH7sWyYjyeuzsEo6YAKjYkQvgEIkknU7Y1lhfwyBvGeEGqg6RUcKGoLNXrWMNQ3PKQ
0Zh5ZE594F/9Fg4jd9QcwM/aUimyQCGbgvv6q1mzbbwzjMailSW6603y7D78WNyXtzchTraBlHqe
vBSJXA9VaEKCUZfXekuW003McJL/7d4f8dbz6rmNBbf1C8OcNYawPwQ1yKgYnbHWrpf6M1PQ3ZYZ
r0dWW/F9UG2KJ9J6unPxyrz5w4Piwuqa9fNkbCYF5GELPUY3M0xoB4ql6JAGYBHCiiTWL/7NkPlD
3xFo89m8fZhe34T5TWaqnoKd3AS+J+LYbYXY2/AaJEQ4kMBGBjL9y/tS3ia+4BX9Dkm0bz+51u+H
KMvG7CZ/mblBPhtHtrqqMSfPWpl/tfFAxEYgDsk5zh25JvuOmapnY2Qf93BL1O/BOuiy2xnjNeNM
kUEIjAtIt3/QsC0SGSes49IQlbn/xGPNCwIozxcOFGoKANAmCAwiXRIRc9XNfYhXNDBOIbb4mnu5
T8khnm6ZHgBpUEFOHHbz49WZ2TCUlsp4VKROLFEYiX8BNERlBUoca1PXXi9kVfmNYPjaCfMEFnI6
XH5yaZGcssSg9kOEirSTf6AyyedCP+u7kRt5j1jyjBusp8rjhs2oCmNB2SyPQQgHJwH8C+R9FP2c
GSVKUStlo60s1RNVO24CyW1DXt45WYr+j2A0yIn8qWoobARhTrcLrfiABSahc1b6TGKsGngx6kD5
EH5YyxRj7FSEeCby0iB8tO+WisIoDCOoR1sRkBvfIokUc1AiILEksh6Zvaa+ErzuEbTHpLAlhQAS
zhmGPRO6g4N2Kwz2rr6nLUPtGaGa+fyNwmDgAvDgA7oEU5FsJL/3cKHcuaU0V5ScDxKsRUCQbkrN
WynSnkpfD5PYqHrgINEbH1YTn7ZQL4DL1fsLG9xV7/r/+tR+xgcIftbeKgx/wzxHWR81JDnFid15
oJMlfWW6zYFkXb2Z3YQ/Z4MvrA7Ogj6Iw3nhyxQs0iwTnIhIJ6WMqOnqdPTM4yj9moaln0vrXwNX
hLW3ZLoW1Tl2PBFEesQuhLfbd/Xhv8BNQ0Wpa3N2PFOlowsAY9cgKbcvoBFLZaA5RN9rZfAHpTI7
BaUwOHL923Yj8ioZ3Bi1BQ1641AoFA+GWqj2IXeEOr/mI5qAH+t/g0rualvIF0kajyGbtqsguBOZ
hLFJOrhCsze3xPs9P3kvi8z800IsiLr8BfLdpwnpGGQ4znMRFgpaJQsBBQC2W4njVkuRIMU1j+oy
c0R8Id1pGnurnSLUqNjOVBqBPQG3Cez7Cb72+vtyViWjIXuOo2nYe/sGNqWKb9jj8Ipr62ILL6Eq
lEnZdPq6571hwjiM7ZIkg395w7m47eReyntMmIXznh3PTrv4W0Wf3WbuNbyMnR0HsZXRUZxytILv
K1dXow2RMqWbrbqLoR7k8f1oyeW61PwrigXa3GejLiILM+VA7najCgQB8S2J/lp6i5xho09ZcWfk
QjqED9L+18RpirlQ3i+Gi30POFoFjQYWOjTfQDTsE5G/Pv4rWP/34vaOxOCfedjQBzPABb4wdVUo
W5B7ch+YFslfp4gu/sqlX6ffM/0JdEK9pMhNo2pFjwiVJZ2dGczL66FqAMg36ycctBo3p3tkMIfv
/b8SxE/HxHKfP1lhee891e22UaaOuE5ydeFzc7eM1ShgX3d7G2Fj6DwwrIF/mzqqbjhU3Zm/oGzX
GbkBOVNvE344/L5zbFfKiLFUalrhd7LfJgGK+ng8nZoXA/WE1Yt+gWSqut5M9B6Iu/NBsUV4w/jz
LWclFwwbqZ267WPLxRhSb1aVCEucdFGh5zz67iamG4Qc020w7huoiqeynakuGMYadQJ5mVcf5GFJ
ZWME6tFkXKkzl3jsdKbNeaJCGe3iE6F1Xtr3x98OHZtHDZrUPar1qBgpccveASam+bMo53sFnzZJ
dzakuUlfhn/Pzn3j0QxYFxPNMo45q4rcpBHILnPCfv0xygUtdrO/oovkxFUcgY+yeRAwc9tVGlYg
DB2lKLL8G8KUmmBGyecE0gabh9lipZhuKMrAIVUprNtAlquC5jl14Ihs9IHroF4USUZzd61T52R0
Mgvc7tRWkFGtXjZyHtXp5VD7NSETyv1FUqXnEn9i4HreF0pyuT0n0bdgqll1D8FEYCf+GG2TzBjy
gNH6rgF3wYXgpFmUa+6Pw2RjFIeVWANUoCTe4UI9fOI7H9WHGs0ZOqQDFA/MZI6hi4P5sVUU94fh
tHD6YoYDnJlZ1jSeWg8jj6iBVtsRNyQY6qHnOIn/2Wf9T3CfuGQYj2niEs0TAeL8NWqculBpEWMX
YHHzCCKICID7sPD6SASLkez6ieMTsEZnCMtMHRJNGvRoc7anblZhmXHIwE6xVRLvIJEf27MRSEBL
kVnw/9dIlMBQWoclI+IDFwLM1fmNWUxMyg7MnnTnCSDR8u73ox+aK8b2G7ZWBmVX32thOGslF6mO
DPqqjeeJzxwQa1tVrJYla841ERNKkPUlf/wL+CnZ+Ziyek0WVExZeMHmHkGz7N9QV28Ca90ioDcC
SaG3xXhC/lneQlJEdB/nFc8oiH5m8eXzthwwzNApFzCC4hjtIYI9hUiWKkkII2ieIrqbdoiG+X8f
VrW+fw8qjzdCeF6QoMpItQIV900xZz0ZZJv57545VCOVrv/kNvUmyy6Wb3jD7xRwznb23FHM0a7z
a+wIPHI+HJmgTLWbSp6iwIgx9viufUU7SK3drLzdzlonAjQi+6rf6lvWghtDSEyElYS0e4CJzowV
QgRuBkkxMhQOifipboZ37gdLagotIaEFfvnQPX4WpFUSCRop89xUuHW+hubBlAn3beTzIYVdsWu1
pJvGy6fKP3H1zKajJRIfVu0tuleOYJu0TYYZaldZPC3RRafrIW+GBNFxxTZEqjRd4EdXGCgCyxlo
0xcjuf1EPNyK6Na1mUylaOLS43oso8ixzwrRO/nDR3GmVcppIe2ZLiEMxexpPxjqrbL+Oswpj2iy
3Iil4yEIO5ajVaJtyyjpUQpXtAiOnoXYZcUDFvXDQIE72Mgz9lC66omwWXsaragnd6n8sI81wW4T
kbAF4RMIPNyGpbIHDgv4A07vZtcD1Otfadw0TLuTUNPLwdUtTlGHQ7kYXHOiZYf2m0NQNgfceJXB
CSMFw6PJiQcYMVx+ExcvPDknR/bXEJd2yZwbMZA4q7Sc1hMi0a8ZBCfaUB0NI9cJZDZ+UXnYVt0H
HRoxd2EGZ3U8cjUTSigMGqE5iqJtwDpLUSTwgoWNqbP+xZVwgyHJAkNdxm3+yOy9QpcnfU22JyYZ
pWPE52LxhqUbWdB22zfrsqtkRrUQDQLBGLsDihaMcz3J3rccW7xZQqzDGOEY/SLD6gloPXmIZfbq
cJAO2ZKHO/AWXn6lCNKEOZIpeJAAMa1+oRp/xkwREh55jw6TAlwJlx3Q462nEnonwIg/BbFXZ1X7
+RW5+rWUq6mQQy2rEJF8so6nTJxSwDnmimLWjcq7TVHOxtphJKmJPQ4DCd+zu98ao3jQnq9oKZen
/mdo1xRgAQQXKzy983u+Frecm+YGXyGlc0tPAvf2V/jg6HLm0qfYPV6zmTx+x89b8fn4gaHE/2kV
tGKbHUmErbsIbs+5j4thGMb5sGiNzBYkvHUFFXdnJNvVoLUFEL6J3sJl59BjHvPp71XfARnvFSvm
eXp4PBD7R+jl7Lipas9BwCBd2s6sX6/5k4lDTaVZ3D/0513OhlVHxK5loIzAwQEpOjEsRSAaZk0S
uvB6KRTXnjqhBCsNjN09wlEBtOpvjxbRCtMhs3ALB7+cgruDSHHbn407ONwzY0j7BNakmujmz+Dd
fDwOZ1Uk/tvfkn9f/jCKNuOKRIWD+RO7kKeWjR1OyfzTQ0ULC50p8n3Itm9pZhjYV+1hOLKDbXnP
iAheVUOl9Jx4lcbog3s4Cv1I9BGdYO4V3FbXy7x9LmQGgQUAmEayfSnFkiWxdxQ/+PdIsuw1GDoY
XLwdn1SOr43aOBXuV9as2qJ57WjSoz123SDszrW/KJYSOkBgQL77Fx5K8RLuSJQp9/mgryqlO+ZU
ayY5rWC+jd+cWNHCPbrf4jv8Z6f/wYo6SK70y+QK184m/zrQAnx/RAAbt1M1y1fXdcM+hUzff/Tj
iWCE6ngm96Cib/bsCt4nVP1C1Ma1JEtO+XZMyXdhO5JH8m+ZgGbzR2OYvzaxcSmIWuXDpERCOpxN
VIfxHwjb8nlElN8LWyXMYblDXfvDCqZJmAmu76Vq/MbMla0P/oPqXptybyAK4EZnSVv/+y8jVTgD
aWLu7QcxFD9fN9oowyCGH0sTbUm0xC7uLu5Xzj2SCqB1EjR0ujtqtkcxN6OiTsdQyfu8PXbgc7W1
YXommgNMbXeLu2xHqTnrpTwL9fT86Qm/ntfAIUMngrqxKrDkGbhVsfXSJlJQg7FmEfHh6d27pw8b
aGbOhGsGqrdAJCLT/o5Mbjvgp3KtAgbWRJflVrLbf7wRZqrnHhNTX/ljiLD1n8ocMmSRW6NukrAO
OTXJq5Nwd/C2P0Ey2tMIMKSUphkhqDSfc7i/Et5QZkO/6UpJ4nKrKc/dnBDmZ7/8njZERxHpA+CB
vfjD2Nd3Wj91B+fWJt5hpWGy8rjJQCIeJ8jkwpv5PzNN2aSKdDNkBaW9Tg4dl/PA8qmyiCYarrDW
ePUCJ+/AD+L3p///ScSFMPQ4N2QTsdqjfOsgckv7jsuZEB9/eRR3RcsZHHOn5SAjZmZed70Q2Xdl
pUE5jXWkdHh45VEiKcVWMhnWvfhnQWb0VnTTi47qsr1661Lt0nQ1otGCC+4YvdOz73QHaOFjqTuC
pF0/qiX0I9UWAEW+SZfdkCuYX8PWYIJcY/nrc6xLD3s05iJf7luyejynyEeJIew3akQUl6tTwI1S
5lvzyWJicqE8sVOwbopOkAaC8M32KSsT3j5C4sZ6ZR1HiA7rvgw6oR7CiiQZ1E9N5F25t3cZtG/8
+Prq0a+sYZqfoSNOOX9LGWmC5ppynV4xuy9benHdYy5aYrGIK1kbi7WUZv+ZAU8t+X86hnt6NNMU
9He2NEg2bZ7abZBsWr2w53Uv6ijRkJvlOAQltW/TQg9L6D2T7pLJeSefPTNS/o4rc9m0Qsb/RzWR
+xfZrGJOYr2+c3PB/wHh7OcJeRvTS6N2rAdI1QQ382/Vn+TC+NmRNezUp6TB/KjnAa566N9oqqPp
JLlmhiGoey5BkMD+0E4azY1caYVbRjmlK5X7++cAmGc9S/kqgkoNegR0azTqnls3Ot52U9qL0V8D
t8B4dipb2qwJTpyK0tEcqEkTh7MdLECmTKGquG/vJpd98jusWsrYAE2r2o1N3uHw7xJ9ja9cuw1s
qUYLV+cpFt3NXnU3wlhX0sMsqDLRts8/8XWt/mUA9Ew8Qfwn7kmmbfNbQ3845tM4MBkGmCCRkwuH
AOH93nUAzwc+JBWtfsO19y1xErpGCu4XXR1HzGWvxjhCjFxySroaFJkWtaDABy+1zvrfYEtaFkVH
TX535QpjHIVVsjhC/DbJRR58TsvEQZxFwb8HlWwSdVNbLmVyPqtTS8a1p6De1bfCuU69FGwgTcoC
99ego0DbIYtxxkt+HEZ1g2lSOL2jV/p5zqP1F9HzPSQ8DiK5scfk15aZJKHpLShdUpkxtflCQUC5
mCl5Ho+7PtbMhyob5su3dF7pODA3wROX5UdzFls5ju3/e8/PQwvJ2CsuGhWnNB2nt9uDT7cBB2i3
wAhYnBWODdACSkEpAlol1/maA0DYaLD+tX3FPyLZrBQcpNbaR755nE6DJnzN0iB/UsqjJ1Xy4iuR
461SZa4HKAZyyS8Aw32+JW8BDRlJKYUik5A94SfFxwdURgd+YdN5237LZDMLTZ6TRyWS7/9G43lb
GC0typvjkq4kqq4gTO/TZE6CytA+6EeAA29oFZfQoPxmn0PmLn4HoKk0nhGZbv2MQOFBJbFCWeJ4
WPG+47AlDKHmIOe9lJidSfXMHqYADBSFGTYHRhAEQK4IZEIy+MfxRF1bR9yA2wNKekXTQ0B1586d
z/r8m0vNtft0ILpUMC3uVULJGVMQJkXy9GIlbPMQiD+O4KQPnkpCWH+Lw9d/ZmHV2LW7fzz+Rl+H
/D4NHn/ZFLsO7U++3TWzj7U67b82q20OKgx5RFsntcIdRn+d4IKZUNNjbsIvGXM+aA9fr/NTaMgS
YRZISDyZM5RTTd3ZbkBsrfTjukFllgpzaf9Ome61Kry2RVbFBm8pdnzCXmYVDzUmBn8Nu4lqLRhE
1PuVYUR5fjxtmjS339J4ApFHDMuU6YrVwlLy71gGiqydxq1j3jLDoHVMce+ytumPKu8am8DaG+xG
Xm1Ts51p9JWdFEm4Rz1OW1uq8LaVZ/h5pENICL/jhp3ad9knTITlC71Dx1C7xom0OZz1SQDz67Pf
NkyB6MCaDkzpnggGvB3Amsg6+lQb4jOojp0eo9UYNhCEZ/Smr/LRPigXjRSL0G8hFdWVOM6I1w7k
G2rj23Vx64YniALICgCOWcBZpjiHiFR8YgezBzw4o9usw7KyZwSUdAEqhsYEeKStsYkoGgpRlO5L
n5gQMqNV4Bb91QMd9WTl/uZIqJbpXINTDxffBtahH90DUnVlkR8/Wsy8b0SEnyqOwuT5dhUp7DC7
C3BAmGynmMGM3nJrfJeNxYSrgM1EZryr4twoQUuIj/WxC7ys8L61f7LSS9Mj4jhFtOd72YfSjVxV
tsYFp+Bif8bfKJz0ymtLv1tM9SuYnFZYYDrqUlFu1QR/g9d32g6qYrl/4BnL5Va5bMBIuIbDOX2T
GsMdvG3H0e5wNbzanVMz3CJnWd1XUnhOML9N0T6PcX9jUUaRpvvwxfv7IOHWwQvwjisWpJHdvFxj
pO+Yb1/xrGmVNprFR2MKfd+GEDAYawLM4hU/0vAGZnftlnwYGLPBmmmLfay3fOO/o1UVjaGcBpJf
USAA1bg9fdaRdPC5YKFS9sYhVP3uLodz98rPFlJqqxlbJda7g1YMXpLfy89H3C9auh78mlOckwMV
nF/qWJy+TCsmM8JANBK7HbcZYLYmwluU8DDTcQwEsqTteoWGjYrAXFYdhljsax/PZZvF1jsq7mpv
Jgi8dldOwKNswlkyas6Tk2ccqg8OQTrkafmVJtxcecJ/6CqHZIYIEw2l3bTkAR6uCz9nB9FE1hen
YHJ6ucKU9derPdDZ5eAih+DrYa31Q+ylrBex5TfCJVuCTh7aPqVSznrNeHuLCAGAiS7Cr7psFjq5
iCmpr2cFRag2PGYdck8Klm+iMTGUjLbGz/YzSW3K887Nvps2AJ0ZYYukjPpo/OPGsYXEzgr528+g
3oJYoYwc3rj2Ya6ZM5K85+eDzlhkU9jOAwer8QtaWXxO+ZN0Mw4GeKRDumv2/fW/jWE4AHTUGfAc
l3Dtvx/KW4rSES8HIbN6i/fTQm3QoRtmJ0lXpckCxFfjIlE7CQE4Vudh3/NWY3Q0Q8hX6YhHFu5w
k0BbfRSxcI68QNbc1LF/Q6RO20YpiIT8xJZyAX8P6YGj/97eRL+dMA7Idh1923/Gz52cAU9ZdqCq
WGQ5BgYJtO+iv8CEKWzybp0hvn1omehDLSjOMAVQ99dFSh3C8InIpAu2PFfXhW88NZFPlYR/Nyyy
w53wnSV4rbY/gdQF8DoXeKgPRGvVBv9k5OLZw00y2zf2WdMabTxb/vvFf1pZA6eSCxDL/JTxsQ+N
Iv59x/cOByozVYqihHPO/6KsGsmDCG+gXxssrnMowCJjgVXMxB3zK7WcWqucREdTj2ufJ4TWbcAx
9w1Rn64J8zXnpHbiJrqNsfdaSe2GTwdMXHliBCBIVkYZlII5Y5SJtPFvbvzk2B2IYVcvo2MXvDmp
qbKWmNA6aRk1bQcvv881kEXZ/Yl/Qs9UCltu8rrNLrnvBJ8odW56+yYwIVdzgwpyrGIV8Tg+v+qt
yK0C6P2fA70wmHhiOvsDqsIj2bLA6JOXIjQh5kOQFuamMfRj2O/vwec4/B1a/fLTv3PWo1L4LFHe
0oM8kzPXv3QJqPA+iWY7Kahe3VRnEl00bvIeF7qeqAQUg8ffRqTeExnzSyPpPhFHSzqE4XlEvJWv
jJc2VCcKA2tLWlZI5EJAQ5GZBJEDP9bJcVhr49nfPXCXljIjHtp1goWR+a39XE5IS2Ela6F8X1rT
L8GLti+GeZ71kGYs0EUc79Q1CLiW8XFvfWANR6bYrcOOA0W7a6xljrVboTMReZKL3ZpGtbtD6Gnc
iZItl1DgoKnSqZDc9tEAiqkS8zFYV4KChmO41ohYS5+vmS3VAFfNi6ygJZlTasN9B0j+KahqifmF
MX4fa/QydXd+X9ectHllJWmI32He/g/H1Hd3keFyePQSNRj9Ex9k6zYW/JLkEw43YsTpa27uNAy5
pumfLJuVfzwZsnQe7mbJIxz2IW4HKIJDqpuyJLTBkwsmc2KM84lDbxCceeyCCV30899PznIR8s3R
HpscXDmQpMyfYD5/ggdEoXrydsiHAz+6wATRzZonEqJyYF3GmxD36Gt2jvvDgC8n0TFb00pLNQI0
XMVr4azUg/5GWygKbUsbR5fly+gIMv4UASM9HC9cFh8oyWAAVVpooXoLktQLJK4ffExSPa83/IRM
dpiDi4sDDZVhZjpBF+5TtvXZ7VW54B5Cd/iyNFbY/HQMokKNr+3FcviFKto3ulhJrO/aOf5r/e9r
uGADjJG5HoFhMlGc2qe/zCON5BGYbfxmq9rrOq4RxMgXGJJh1201c9P97VL3rlygHTN1/+PcfPTg
Ee+6TTyndyNdB8olk8gtoDlqU5lxbp9blMi3C5SNZcw897yoBIGD0kD4mjGQeTeSP+3qWfEmnNG0
YyU4wrL6+IFLpuvqGQ36O9av93kNw+NO5Mx748eCw5ldXAWrIYQKUOFcl01R/il8T6bbz6qYiuKX
jT0aDl5ENUES6vcBq8+74VAK3nV8/ZfAwyodmaQL0+OA7Cv1853AnY9LmosP7hFIEOk0DG5uJ7VR
kXgon6KyZwm3RUfDoatp54eC/aE2QDchhMgCgce6tUfPJ3m+n4jcHg0UUF6N4s6cuglK5/cJ9Z2y
fiJW8X8UJ5eURy7t3+qZ8aeCow6bqcTRR5qvOX+iL4dettRykIZXOCON/3g0uzQpBrTqgKKvIb+e
1FgFf/vsIJaKe6OYrpJv49KWB6GNniMIyyb0T2ZbTO0Y8z42oddW3Y/HIRmJdxPpT3mcMxh1rFvD
gzwOkhfYosojp/bu34p3JAXGmKf0xHkT5IkbYtMmR2jOhgyHxHUTRr8D0JOHFWTQl2NRcxQOexM8
scrw1mP/WCmTnlGby6f9aSBFaCk/t4KjO0JVKjnds/5bcLB/oJtcJtHVCS0exz6vQhNryY4QJhrW
Cylfj3yAjcag4axN1X3LYKI/STaAKZM+JmOMwCtkFg70ces00f4zDlJAa6WLKBzaY18p5vmxGAcv
hvhGT7HOwTddVpM9odfDF5M/r01ko+V1LnMVeHpbNeBv1cJjX6hUNSKCZlJ70QYcS6ZHOYDNcc1D
o8y3zCtY0tvpMXj46kJsXND1xnBbFJstguZZN5DUrIBU5ar9x+z1VmOAFg6X6oVs/MZ6YgcWkuwl
BNh/h/fRlwLwdF+tvRGUySUB7633/fgi4dedjK/z+UoW6LW6iKzQfMTpWJw5o5ctii5ixLZlqSI4
SidIzYQiVx0aoHArOySvLC//3Vatq+h9F/jgX09dlAX+SY+fyU/X7LCZnTsXvWSM1cnDYu9XD8YH
xNKiWL6LgxJOwztklnsKzePn1cPowP+PG8gLmU1XoOIKfGtwgOaZIA0NvgzduUM5hNtgFDOSIB3d
pAmxTL6nx4Htldb8WE7xOlf7jFlmX142SZxJpdImLsMxpBna5/5l4Wgyxe514p7YsQzxFtMvFAYT
l1fuEx/CbcequGD0N66RfuptG3s+VwRDDeI8kHFc+fd50/o/rgU+G82zAaClS3SYzutf8KGE7yQl
KLQWnPbXK+166U1lz7lLdrY+NsyquYc4HcjOcUl3fwXTUHzaqRuTXXdJ+MIK47kMvU3aaoFWvH3G
hH7jQaWt+JyGmqncgl3XYt4NTFVqbtZZZFjUBz0Bf/ci0UvzhH3UjIMhVILIsDOFOiU6lA/TSgik
+7EDEJdaQVkk7gRbSN4+DTke3ru6YkM3MDoX8Lw9nM1yHZ2YMueS7fYzhabZbKh5tLgK6HHFJFqC
KwIy3AkOEJ6kTGw7VUUZVFfNJKUle2XbVMala7lT0805zKmPThNTDnjlNRmPTP1bZH4zmsWRxkJn
cDIxzD0RSszAhHZOHRXE9o5dgZU/OYMqI8n6rtFj3/73T0NgfwIgckn7EoCDGL3IfTnFOAGWulBD
PZnn4VIlIfcMWusxuNdaSRNQxAnjj3zRyd8IraxS+1xTRiuX/7F6H9Qc9LLVbAHUwN+dkGrCpfHg
J/0GZmUX+AhI5nZ49r3bBOIPFeWFhyn5QCfmb9Wupg43puTld4kXk+Z/4SdxBQSnTb4TWZghxPx/
HdDv/GioqZ26jHNxavHDDjpY+W+Kl2fvOqa4AA94MXicIAlQe0h171WYo/th5PMElaePw2s62Qtg
DOQHw3AhQoRLkgd2nGdWkbQJ8ipdjfw9tBzRQD8aK+qjPrCWq5NJWQ99SkZWux5bE9BMz3oIElxY
cH0x36GabA88Lspu1PFxgrWMFb0zaAf1m/8B5t5lhsgignQtb0G9B+LP6nVOJCs2ScnFnYAXTx7x
8OKIHyUVnehWbZUm3IU/Yb6O+8WtSME9XfCKAQjFmtEGcqkC5SKJCq8a7AL2qb0qbqA7rf6zWLcR
A8oRgRQlQxSdfKjpODglcbfymJUpWCsJEHpmmWU2PsEI23m2XzLu+ApP/5cQgTs7MrrrdSCBpnT3
DRvIA60Wn8eMhoLO79O13UReV0/76IbnD3ty01DAAPPbXnBpay/bCzgMIqsEEyPN6Owivym3NzzI
hdqstvLADG0zqV1u7WIUyw2ZDEPvGEtSSypVcJE2bSMXbXUJClC20xgZ/pr0jafZt0cbHfMRySiH
t3UynoiJB0Tvng0ehaoo5DDk1mldLOOu9Uz3ysB8uBwtEving5wZevNt0phVJbjdbiMo1sDyi8zW
f7PCd4LTnqdo2ByoKfX/UPsoW4aPdjbV+Mzf53I9IinOkJKNJdjjYgqgk2nO3IPm1OhhQhJhy1Ft
sVAmxqyZBUKOycdSZu5eYfEjFQm7kbj+YB4DQ4zeFsdTOtxMcx3pgTe140MvflrPDbq1AJqIhKZ4
Bv0CUUuMwvtH0sEkl3aOgf0SX8fMAjgLE5ynhH60fb8QX2H88KS11OZH36v7opUACLAcOftHjoRK
zaACm5hkHzbzqWLAfAOM/e047ab0u6VXYY14PnLHndwP2MSQeDearg5/YH5iTVSKouwmhjUStVgf
THnf4EyKtk+SOtcWwsl5e5CCGQlKkMxLmo7mSAHpONEPPGcvEDrcrLFa9O6ZiKnUrNMomYplkyqI
eFmzG4dAgQS4KwxetjDhyjYR3tqsalhuW9BlABCniyWwtEe43wvwX01N/+iF02h0H+y2UseNds6V
iD3sdeuglsDV38zHApbBKHYf3mHyWI5k2mDaaPQATyxqL9NlmNuoLvZPEFRpn6Gh6sf+bsNC1zMl
h4om/SCdsqh5F+I3mBBXNfLaA9ZLs1YgXNdCiyxKwH1qTBZwfEnSd4NWy1bJxgdPVOXzCwkI37NC
R4Y9eldEdbvV1Gv3mf08Gl8dHN9s6V54XKA+DHLa+NG7wMMtRMZ/ecTzUwNkXoNPVKcpTD+tJ+Se
rmHFlpKvdYo93J7iDsEpiFkeeTJPMBiMglV2MzVcAaxnomSlXQg2BfHXD1Ny1aAz5tQ0+wtnZ9hT
TTzzhd36TajcQK0nA8w72kXJiW1F/lFWV5jW0vjVOz9UAFgFshRwq0jeI6xIZpv98YzwOCX4MizM
91wa0cXAReQMcmHNO4kKNP2YzsYl1ESycTv9KmjMSnmxZbTvt1mJL0Zyx+PTeUEpPZ4ijN7kh3yc
YzvStxCmwgVDrQcWypDkJ16ZCftembOKhEducJRDWOB/f+febfktK+j5UwTHUblCI8WNYetG2DuO
fvqCFCzQzuvlSbBZNEji/4CFKzRT4htTqo2LxYv/oRq//CyND8OTRsktTJ6MKexu1PNAww5hYeki
yEmM0gzhWLwtmKC9YlJ2WoUFjUJxLl9BlXSqc/wi6BmxtnSqfcIruPm7uoYImAnoaRzckp3/AGRp
Detaw2jKaM68Q6az2BNbyT2PGciR+RkdC63GqIlhuY6SC429gqe0XVXLEZQ28c7ZC1uSBXupvH7B
0rAsLMe5zj8VKeQNCuZKIQlDjFqZGDmpi6OwgVUeO8lZeOx2m8Z+Jqxr/wU4a6O1BpOvlEWtR7a6
8hMAUT+M21HBZGg/1attanEIKRr32xLuHq0iTgVN4SpUkddziLXcGD8MYZz/lRjIlhI4DlUFcNet
srMjZ6SfYP9D4mc7ZDDP4Ha1B7m8j1rDlu4Ht2yEBG7+1ibp1HZCjQbJrCVA5qkGxtVS1qNtTvGN
mnFJLm4ADgVpka5hatG1/JhcFc2y3KYWytHpGy4DWtt0WKOhlfclPUj0cHL7ByLBDl/vlkHxQ5Zr
r6yhgraH5j896G9EjIXFyUU7smlXf76vm1AAeCg8YWPS1ZqwDUIeztez28I26IT2Fbyc1eIOzMQy
MyIlDNkh4NOWkuq9YbyxspRNE/F0FfFmM0ZkX4FjxL2znurlM4Ub2TcQ5ruX90Eh2WvxMsdgliLf
38/+B1iWT2HKTp0yfMZPKDbtEMoz7gsOR5DHFHt4GUPgAjsOson47i/N328SM+MmrfOFAdzH1q1h
xRhrTTKuOqsWh4w/sD7oJQTySvvQ07wvt0Kl6RTZCeJ+BWJ/aOxSiX3q+mq2w6NtzlOaqoGrO8GY
QVSmg7eCt/sVs4M0ebyNvi8dBf4DcD4A5MsFicIVY6uHDy0ELK0uH8kUhdYh9fHWiH3lHILlPIDg
7Rl4k/Rpj/eWJCo30lCYdBUSiZpgCLTcYo34MXuicGR3DpZJ9QpX+Nc3VXiGpluDchwCBNZumjnr
dss3Idr0lggJ1ZlJNCTaKSPHhGc/+FenCUPfHNLLDhV5uh755QM1WA0zjVBaYEYbiJqh8JRM+QFr
KqW9/KqZMqfr6z7bG2lUE/DakVfXUfMzuhg29yKa/ifchgcsFV+16EX3XZ15evL+TnK3euAmY6Xg
NEOFKiWBW0Lgg0IENuakiiLq7hDiytxFBUcKnjtuScCFvX8pI1L75zFQEyYxE7D0C+vsGmO+4B7C
JNtiLW7PYXZqKaeYCySsnNtzmsNNAUQrC3DzJ2hXgiNi2F1K4k3zfdkVriTkGNJwc2GlY6121ENb
dDtQRIdbhLaRhJU9fyOo72q0ftDan6B2Egcga0ToITEJojnhiB43KLZV6wxvpLThrPCFv/EGNq4z
bBcOq8UUT9FJWj/PRsUI51btiJW9Ro5RXPLR8dGfLuI30PnYQcsBq+nuwOEA1SHwPQ9utDDfrJGx
PzRBnW2Qt64Qz8HtB5bsT0UfwV/EiXoMgdQPYEI28Z+GcMp3n/6vJUVL3vxX6k/yGkAPPMjtETNn
0NeB/XG80RyAUgxOMwOQAigga6WUAV3hA4c4EOYuyLVO80w+NrZIWBzOXCSSQLrZGrAh16VuN9OV
t+k2HzMnWiZgDid8vWIkCgJh7cKlCNW6kK/cd0wwvxMshhvujOdENKerqgRqG1fBhk2TNfLAFwsg
ymW5vzPVXS7j6q7i4OzX1gf9aoPlpqXuunD24xlocYg93qHipr/ui5x8KLi+x20bgS699myjEemb
nZrdAqTLEtzQZLUqtxnkMhpmFTfKI98Rlz9+ullwi8cyedJtR/3mA9HYSL50uDC40zctqlS3CF8G
BWliJka5Lo7j4hCu9a4d0dDlmg52KKGxPBm//mOl1lSyoZjf21D/NIA5FLXPNKH4g4qcLB9osgwD
+jurI67cSYQLubgERl5GNPc+4DsWCzvcVapoPkuiz/8mdG+LG85ZFQnEYYYAmRJtIKTwvZV15DWn
uy3LgyU6KNwHpdrBHdiivKvls8JBt1Ydsj5W1KfSzAbU8cDRiJB2uNw/D80j8KQ1BEsQhQta6LsZ
9OapVVTIvoC/GmYpMpT9GcI6hl/sXyKUKz29BjRCEuJq1M3cdjVVbRCu6F3Oaam9Pv5eChXyLeZA
NsUVWK2a3X6TRJ/PUBybsBSOWVgBvEFulnfqfgXDCkDndrj78F1FnnnIFcov+4ebVOKbxEF9h5H6
J5wTKYqY4bZpmauaalHkIh/XB/iebO43uTOxdM02SVGF+xVUiG9vDcT4lGr5Vvp0R1Y0hoXPSGNi
lFrUNMty9tiYyG8j1Rq5GBP9ZHUiWigAVsCh46HBCK30D7Ae46ik+6BFz1IPkiCXk+j13ctGP6HN
4KePdnOc0AVLP2RtzB+80pUJetVJpyMhVEB196SJcscStvmX//8MhWB+VSyR+CtYRENbrEfjE/4E
TPABYe3XWvzTpDvg8D+DQVitPm0V4170hmIwc8Y3yOpwFkOxAdSMVK6Y8sEv8MH8S4K2LsBD1A6z
ceoZWyFu+j8z2ndjfLp6dEXFjQuSthJl0Xqsy7DPvyxqmlYwmr7JuSTRVFuP37ZPoKWXRGD0EI4b
Be/2HxbpAz//45mcJaWnVPu44p27n/OgXNvOEW3Skj2rfCdLA8bfCmy8TI8dMK8TZyFyd7fFkjxI
pGCsk+yJ/CsJEthNkYDvdaZ8TrvLhJFP/2RQIInLYrQwerexD71g7dI4f0ts4oJpr643ErPu9/ia
vNIHzIpWShq6kcBGMntDUzCpoOpT/bNwCAJsiopwYlWxWk08mwVgg9kYEKNtXf4+iy3jKsgjSDRg
dZ17J8cwM8ZZYPZRis1qwzr/SfdJFdXWnQSOpbHUnYWgapfxsEq79qmEcqCJSWeDZ4w5IGY8O3Gy
zfIOVf+hvCz3WPuM+ZraCNyeODBem/p9dnrx6tNP2Rt2umk76dA94zIwdc1ATbWNGSybEJpONjUU
MIr9ckNMuU6MJ1lLMLvKvsD4kS/Wmru8Wz2AOdsR6xPvcl0GKS+bvfiCWWPIOu6RZRm5el7O1T7J
FvEyLxYM8q+18iNIyEehOSIVEqOgdbZ7wyfWiqO9HTkrf64QiGfjAiRMRYrPcJTT3yzi8PdGVAqA
i+TzAjW9xAx+iApb8MxiPmU/0LmffayajRk3d+GT/CJUw8XMrdllcwuJpLSg8Vlq6mbWQgZhVbUs
73eUe9XUcj4yVz/d+vxfX+AznmtOBK6nY8Ksu+312gE4hsamvXz/BDCExMnOjVC5gXOdrRSBuqyf
fUEBc5AZmrzcTIDML8Xo5PLN/Zopl3N+CE1ezFL0JefxThyw8Ef/NgFm9RMMEsV9wh6xNDkAeTjT
DlX8d7rZO1v4ySmOYv3toxmVUjlm0cQywQX8Td6xXrBiSOyUdjwUcdYIoUX7ooW01OMjWMZNGJ7n
bMyNXbcEiUuVj752BsuO7xN510hicm34gKs/dvrXQkqTBl8JlbjPt1AVgip/wG+FtnC8WkUOeIEK
v1NLv7XPJgCaFfC+KysrjRTFAT7D+r5vzKd9Hqnv3TOHstovCCV8+jEjbRLHGhQQbw44OgnV8XWH
ccmZmWX+iP6qYZHKwS7p3VNLuS2fYqQUSaQcFayY5mY5ZOQ2Eg+qdSXdCwwUD+Axy3My+SQZX5D+
FRX8Z/QOvW2QBeBhndY+wG9Qh1aOcPA/pKGXjUPLREMxgWVEdHPC6vYbHRXv4HxPya7D0aqkDLuS
gkvPkVddkbshETlBMVWAHj/x7bZVzkRhF5snTWSI9OvXZT9Ym26IYAaioP3Q62JU0ExTxvrujlM0
1cW8M9HC/HkeP/ZVVkQ37j8Q7Zt5yHziaQX18NqfVyGA1NRvJ+fR91kjldu9jHD8DLlV5nvcekik
uC4TPsEMpoEoPcM1BpZGwnoI5bO88Yh0rUEZJFd9cwhghzLS4wXIlmtPgY3/eclnEyXzWNtPJaUx
AdC9gjn0M1kcEPcRycvpyonJtPM9+D6IiTc+debVqVL2lxHxKxagTJzFqAw3IH2LlIVL4mxrEmjJ
P5Tdrhh5fQmFJsch2B+K1as6Dw5vJ38WtbnLLx56zOn8nJatm/KT5o+4p8P9jIdJEzXx81dceD9i
k0KurPw817Jj6T5CawsGINvi+0HerxGKcn+oxy5oEZJSfPqNFj5uqhO+xXQVUGROtN8zpjFFDNrH
H9qimRzZHPiqiVhG2Xh6hAwSMjspgLXl6pMsvvnBl6ohEFFy0wPNsTWbnlaIO2eY3hKskA4KBrlY
ABiU3ygsDVdqI/aQ9n6H2FE6IFNo/GjEN+Xge8wdAxe1DFSBE38Q/hnod9b8kOyMzAdN6Sa4J2KZ
r19uiRTAiUuUWRRCVWkaGM6QqvLOaPzJvOMChPu79AARd34OD5LWHj7m7aUNLCZyA0Cy7tEHskMI
XQ7+0E8lMWsckYmvJZqiGMZUUuZQ3V17/qiRxQD7Vj/bOun6dFPcLUeh+NzZNhEs1haA3joyBwVW
+xd392N7lXChkqvgkAZa6zWBrmRr5ym/wyKvyX52ZgPIG5GijkcAOPNhqMPDSuPTXcZuCq527Gf7
QN1M/PTqgYq+ahJCI7DXA+4Q2GrkrvuuXSJGvo8CP+jQeHcPmJvByBYM7TbgC0QqU+OQtUInmAQ4
qR2V9iG8ZOC6ufwmr65IIDfjF7xd/K/dCws480HY38idnBfOVUpRHEbVMYAupLMqb+q1y4Bzrouy
+zsq7z4667/a8IodgT6t2cUpNI3KM5xotbYHCgnuz4+4nuc0InkGG7VMt9L0HZmnk//Tw6dot2iP
5AcFdfvLyG4ruBfrGtZYReJUWTezEMAa+D92E5DFKHLQhX/Gd7I7JTtp8YriLOJuGKUSv5cZWr38
jzC15Xip8XfK4aX0X0JuDNTMy6wOLlG4B50Ec0KWU+2c94CKsSexAK7E42oNxU5Bt3HZ7TauxJwB
7+nbRR/gG6wBX70XNrz+JW4AbyTuGraQ4azhxa3QBc+3m/kKRGKCg9uZQI5Ot2Mv7wPOfYluTFWT
BGJhzf+2iLwJZqpJIhLhzFCtUidU/l3pLpFm/VeucLsUhgPAWj2R4l4oBBLexcVHN4nAwBX1IwNx
9oQ9bZjOjlTIcRWszDGpYRuAuqTCRaTwsV2qrpCnfZgmJvUoPdDKP4cNHrPnE7WBksT4WHeon7Fl
44MongzbPecfZs0PtbspqjeFlf9O8UBL9wrUqO8mmlpdmvQm02PSFEvbjoRKiUDHFtmYE9E2dEhD
XQ+cWULvhRY67MeAWP6WyP9QgcmubMVmw+PsjkZcioT81b40yES1Hwd4ECfkP0xglOjMqkTUtM89
c7ZvWsMAmbC0F5/LBnS0ii6D7l32mBk9JfwyuFLebl5kBzO1IVDTk3cG1E465D3bInvLJBjcfUzg
l7UaLIkD2is59FnmweHNAES+QlkLtB+qTizwoTPwApKJvHT3f+LN42cRVvmTaRL1R60TKU2jc+SZ
m+OiWswIxrGSE07clYA3/1U4p1BzTfraCXubLb6vyhumVpA/7w3sEZZ0ZdGw6QLFGwvolVlKBURa
f7MxLDUCxj9d2GKAC3jEEt8vaM4S4Y8Q2NndK81MYsNCxxRDwqEjVeriUIeK2mhR3aiQ/IjmStFS
hOqC/GI6NJjgw52tFCbsGVfxsuApCJdrpLG8ri0XK2jLFRdpxaqgmUOpwV89ro1rz1lOQSXmf12l
U4QxFFIRtKeAAYn98s82YSRRIFY28w0bF5OiyD+zJuIhXAfpahSydidhDlylacjkGdMwvaR04ITv
Gag/E8xzEtgqmkqzPvzMhZl3yV8MnjkfBSR2fo9JANHIsCSBdlXgRMiLP1TERoU6UgQ+XDVoAyDb
IGin05AGpkD6ZONZ/T5XWBSIrV/kBqygVabvwYM+5ZpFt3BUTRDW/5n7SxLl8JLiHv0lFq1hveix
v8Fda3n42XO8+NLJUPh3Zh11w7iQPmu8cJZgmtYlRmqMTn5WTIaRE5rXXNYqzc2gQkXG8D6AbgQ0
AsPoMxx8r+wBEReUeprRAOztzbY9VSjoTL7csXHVlByuQDfKK0U5D+LceQiT9ykRdcDtX9MCHlPJ
XR/L00NpQD+YwqtwaBKjua0oQ/8blBLCsT8qxg/3E6r1MeGiZ4caON8lNgqi1zEypILvdSVP4ACf
OiHUJiPIkOR0hj72BbAr9uIMGZtAv0JlbidVOs8ldifW2zUfaOWrJGy9dYPHSp52xPKuLSFFhcTU
owBQUdDD8ceeo6ncaCooiaFr3BYtrIvkQEh8PduEaZ8817ScQpoApBYu5XIZIiONxrMg6iG1mDG+
kcnCMeNjyYpDfyBoiNANQJ++dfS6EeCwmWLJsVTVmQ+oEM4n0aT0dsor9W7Rhc08cgfRstt2FVFj
kk2h3MJK6oVUrpPYFfrpaak8onLi6hgbVVLMYcqVTFlunLo9Tl3Q7qJpP62gxeDsNR0hZTqZycVo
UJOhv7P9tXn9R3oTp27G1aW4Xllh4jaNSgLr5FBEokskwgEqpYhhVvSzyFsGPdq50WUJMtd1nQbk
re4qW1h6GsfYLzKO9Dm535QFyjcnYEP8dKNqUtFIJeZbbJH3ck9NAM4Rwfgbbs5jZYZMlYP0z62e
LQ8Hjt6PbjBfv5SQO2FoxreOtPIGY65haP6dTV3+ILrozisENf/WnXdEsu6uCN6EtOtv0tNlPPcM
pUsGNgVw8wQK6Zwl8hXPoU9DifYGyQcd2OcXPu3NW51bCyCycrFPZoPpHzLiifK3TNJ/KdfFbC6m
RFHGh46Wr9E/oxFZWs7jZiSTjYw6n54R1ya7x+AwHwqSr/4ps7iWvwuxzmp/MJwGwQ2Zdibetpyc
jdsOsqhRg7/Yj9v73LGe1YCTglKdC3MGCAP9wo8RVf3gu897XpTuhR5duIYBpf9o3qw3Gx4Zh5Tl
a6XytF+BLgqBFXQTr0iW0WuW6ymes+v6gN2BOz0GkIan5IxSzsi9qVK0cKId8Bk+km6rype5wvq2
T2Bo2BH/afv39z01nwRnv1Jegs2EIxQDYyRtkh8NF15Hkp+Qdop0IzqzmadfRIgFRnrGYpcdjkby
e1hk8qrCboroPHuen3m00GH4oLqvEv6PYlA0RGhzHnVlsR8hKt9YHeXDYrC6zMTIqkNNpHDr+qcj
iPM6oXrvUfRCD+YyXyCY7wqU2mHhZRgYlVS9ZRLLdWaPsdjVSdiTGHpXwF3SCRqdNmYgeTI3w3sf
htFMyi32ZmaliS0HgnEiGLi0CXvTGFAOcTqF4RgU3OpXVkqSfbH3syHZcDEyScBZxnH1je0QFYDJ
eyE4LWAgdmvPVzCDN77qt3k6Th78pTnp7k2J2+zeiUhddjIiflYFa7sDVpzVtyRmdtbStJaXmjTJ
DlQDtQIgOKoHYvw08WUxNYtrJsAn8kz2QJeBaAiMpbXfNdrknC2ahfnIl56BroXvZULmOcEdWYUQ
OpXp9yxCdB1PuQp+j6X5VduNjLkbygw0lnxsH9343Jtn6MHXAqd/SramStab8KrG5L0ZN2NfS7MN
sxToGenX5rP5DGG3yVVV0vASCab/Y8t0QJPkzJ+l7swL509Ut7x7mVdxwCLFcqUbFx4GqcmusKUA
h9yiCJtfemYXmISJD4lRXHQTTBUCmLQqeWPfI03jheNoCmDLEAGcVoqweKYVRyRUPgDWEXaDXULE
RAYBF+vgXToa0XgLaEHT7IzSIXhL5mgTkqrAMLQnvELU0sDHlWLwq7LD6w4WxiHhhIMeKPKgz30E
xT6i6XDcahwNKoH0QoP1F+pyw+nfnAIiSCDDuAciUgV/eOTYTzveP+ArlqDbomYEwx6lo+IV1WSr
5pxR/79cSxjljMItTK/tYFcNOHPbC9bgGMbFfDJzyRVME2nHKE4zWgVS7omMBhauk+28BtVI14UQ
bvLWUjw8LaQG+iQb18r/VlF7tC9Ka14IhkiRvV7PHjp2L3KcbWh2hM4NCZZ7uiLGbie0Z6M05E58
irwfSl50sMPXI2QoQ2Ov5gG4+NS4iAQWhgf//SCYrkhSu0fbrgX7hI/l7pUFh4KW9MeiCcnm1wr5
B3deRPIM1b1XIno3gHQPEcK7TFNBr+Kv5+ShzaTPgfiHAt7wNyadx1jXph1rwrrX4ewyDoG30qJw
YOH5Gp/V4ZT83Td1UodFGCj5lDWxwBQS5scoW1ADmLAQtvrirJPlTi3UWg0M1DqNVlv0abYOgaog
VHp99hX1E9HXlNYIJ6QXeXH6UTJbYUTjVNvBa9IwwklEBmosLaDIvBHaMvVK4KmVpcFdqJgKxo2v
qw1OfmqOA+OSPieAb9PXTv1NOFIs3TMB2+u7XdjUou1KfvBH2YWuwG2FUE6atL6io0HQxmwG1vXn
uw28r2thQ4qZpabXhCMx/eHlrlP/ZwijmdyolfUkR2S8/6QcW5P7mtUq8Ipn9WcfCcPJr9FnwX1/
d5gMsUV1FrwN43GFu2CDDOzxEsGDvW9xUwXPTwULgmGwWbCWqo69zxdmh05f+DrAKtjsFQlOeBmq
7jOaTFw7EXYMTBXm2DnjrC3vsZ+sUSVwy65MOcefA/XC4NoHhLrPFly2bx3aR3StaqwQ1wDfM6/J
uAi6iNvTfV2iw+NQKo0/Io9Izcf79U7TrEhjbd1tphfVRmpJSVWqwHzlfROt42vOtNEjncAhxPLa
sk9yCQlqKYeqdiGWs+4G7OsiLKVh+cbQHR1rIUYAU3yaAL/k+8s96YcyjXrHEtieA95RWZ3k5gYY
qtvB9vynqgvE5dzlHYbmrUE4QQ7D86abIMtY6Le6RLv4M4+5VBgw+7OiAnD2jU0KYfwwvN1/c8f2
RPlr6rMeNWZzTQyoPCYtmkPPVd6q8JdazoEVVYFQIPT43XvNqlcOZ6OgzurXItcdhTlfZkOmF15E
XkeAf4AcSdu3dZrNjdd7dpU82I/y4XiO7KjZXjwI+vPmTG50qfoMyGK37wFvjh5F6x3gV7Ud64UY
orl20z7lRAuz6CYaHoUKSHbP8Ev1qawBtaf4zuZ+IQqtn8sDeyFnzuob6Omn++MaeJevz8cX8KMv
ZGcQjP7tTBnQxhxPgj1MTJJDRpWk8A1v1iOrfoZ4lD6hM3x5WGImtSxqMrfcLzdGK4oO+rUY2bo3
ynnWDrcsUo7QP7BAzw69xkJA8UEUXv7CSKV54fAONyilZbYwmGOSUuNiOeGIe7c3SJNms9R0ylyR
BDdpfUlzuFAAyx7lwcrrNNd09yqAS9OgthEX9o5yl2IGt+Hya0cqCrdzk8NvWABEVnU1oHbcPZn6
mZDQ6z1YA0X83gY1VZsgKsF0baDCdHFTf0Kz1fGR1I+hMEW/wLRWMMA3AIYg8ITleGJUkEyWT/aD
+ZsPAguUDLL4VZwtmIuXgoZinsaXhXyyrt4ETub53PErQVlxvlY05zmbcGS6GiN9u3Wq0vMkuYgL
Bv3dr4i9qFlZfxJdM0qTlAsn6wfooItGLeWQ/5J7eaTbaIndmKAE2VodSwPI4vQndhy0rG2mlagj
xPUuEhZI6Y7paO26UpYjVsHg+ABgGBEXfg1dvj1DRXS3ZaINzbUw6a9W1GRJVCHJEdPKzozqRsHh
ip+ZmkmFerOHSNi23885N0btaSPGzqABUXU60bvZO2LDheZu0JcoCQ2QlzpHzk7VSyplisiuuLFz
+FKXnhaYHRRyzjW18qMNDlyHj/77vTFJ/0UXjNuphCHQq0vsis9qVSAudpeg7Gldva4TJbvgcwS2
8QKqrPsGBwOAlU8DI5SqVMmMVv1mhxHk6bd40zBa+SnYH+gX/EL70bvcA8pIWEbgFz3sJsLxf8tj
lCHRdPfCBDtBFRLu0ucX4aXquWplBFnexbdhJSV5u2BER/WosEP4JLMOkD+S643w/xW4RD5I62tR
MgVWhJ6zhK1wye2Zy3JUBsVJsBpl9CNPF/c1SdVwmR+ueZax4TPyReIaHX5Ji7iCasJXe0b1ipNR
eFHcgQQHidGm9/uH6TwpFRdFM4an2PjU/PE2LwUhow9eUcNyUF3IqnQp4fFk+v6qHXiLwJgdUBkE
XVEcV+8WGVw/edRCs/ny2X1JePLdD+v5OG6dhS0sBRVvi//+pV/JVjKimz3rV5h07OyyBHeBWObC
4b14zkUXJhAwAkVeP1fl0opGiKLMyDk0PwW44XuT+vKGoT/xoQkgzsF1puGzY+Yt6Kndd7/ptJeM
dtopG+bT3UrQ0V7gINUlRII4GMcVdHgF9Eyaix+NoIT9UeFb+23PqOkK1ZyOzK+XOCH+xJT9otOD
11fx+Ne5WycEJv5i7J6zbI7gaUCsUsbF3IwS3tUOCw+tPhfYnTR4wDiu/YsD9/SqljuDZffMmgih
HYa8g+LTkrdkO02Nc/6Hm9Tx1zrOugVOPM1aodtrwjfpAF9mIWHt/0KrW5DmTiTmpW0c/BgqsL6r
wuPy5taT6bwMq7i4Ln24q34ukEvnh3NcGfvSQBUzmSQrrTcNrTiIHL6j/umCAYJGquqCBudGfiwH
U0Nn4Dree+T3kR49xNWxXbiDHc3eXlSQo5zxJR76Q/ETK1Xpaf2g0hCJAiUsg+FbcrC0Vupsg4pg
R5no++9dS+MErBq8iEzLjbzuOPVVNFkOyZFS7WWkwBMmQVSf5FX8MxJXa6aIoZuotDZFbwIlll12
bgPqkgTkOmwYz0881rPAAnFsGwE0m4B4WQOKBhlwSUMZcAXGBvJWnNVRQK2PbMagL/js9Ks1DGQa
wf7MDyKrT43cwBg2SlmQrP93crNvNMn4kmW2yqOa89XYAG84GhTugO+TVne6rhcQPHhqkUg0x2dH
IGGNbuw23sSbQibpunkzDX0XVTRi8u4iMAyQ9tJMxO9ikD0byY7IjSPJSW4rH5T/iDZBgvXCBtBM
E5ADfGIG0n2jXQ2qpXe7tapxulbm7lsHAK7xmEyd/8aXQdMkJe7+Ty3pffsiRWkw5fcpf7ukWGw1
uJPnA2Wpq9hns6XF3boh/9q35cDIli4lJ/4bynYCDGKVOFPwRzUDUWTOTaBpJc218q+i7uoSwJYu
1xqw3YMJViuhUda5OEeRxCWCyOsbzVvf6yCE4TZYLPi3sFYOWmPkS6zNcODKjc+DiqIrKl4Rxfgt
ImiN+9W6RlUWlOBUoJfy6gwxClX2PsfpH9azzbLprwcd4enauyz5e9zPhDwofCtmUxahbp9qjzjU
29JSpUcExdhKYu38U0/00bS1iiSSDzaMYTvBFKX6wIPqeVlDhbppp2iZVP6BMuDk/ebgaf5ft0My
UJSlIoDWv/gAVtlDeRM1TbtZzDYh+IYT2j8ax5fSc/05NWFZhCblfMxURr+/6OKxuKRABEuth7ec
oxtvnSmkedEAWijSSVsLmrn+ydGhHFislXIiHGOqSQ2qYEfxiVMd4YFnrYyXUJ7naf13DinaYVV4
svs7Ys+64svA4iCmHc3dInPAOURBDByLDD9KpcvB0OnR3oEXKpcjv+oySh11qNmKHvNPmJPUcM0T
TL+tRpAvMrOW1EOqC5wUJ957OhW2DuNNWf61VThvGx+YnJt9n3HQmvZmjJRaVyzhfohLNDEVJa1U
iPYK2ZDqPmJlw6Ybgk2GlEEhrE0WBpeF4hIQomLxBwNX9kfGE+9OukeLYXFQXdQcIPy3x6Ig/I8p
O4tpvViqW8l7RVH3bnwjLBqukM8zre8z+Swra220TFe3EK9L990UIGGapJTuKrXwRdLkwMvbeV2s
hSqkNJt/9sLEKU2FA1lNgVJbCR8i4Ro4RuHD9VWs8VbUE5/Y2IsdkIq6tYx4hIm9evUeGiRK5UAr
85bK/WZWndD9gibGj/qX0qaLPiVeTVLRnQO/K1lNhuWiJoJJa44dG/Ptll6Rok1jiNeLSlEgcEpc
5CCJp8WyjnVW8mCuea73OcZwWIe/qfbDA1guK1v/jfEc1EmbSHyOT8ElCLmLkHEnnfwNcLNoJcpv
sqcSFwMNRX9FoX9mfM9Y1pKHT0nVNTzZzQVUC14QxGibfXztcxxQhFvbAW4db0neWmyIeXT1N6ru
2ieiuAmVTEybfD4WeM/CL4AN3prvqToI2UvSJzm14+ebnkW+jFnqtym7TY9ui4PW9urxn26DxkOw
JUOZVcJumCDzKn4NyUnA6KCF5RZCem+TdHgNspyLH1L7vtpQ8DIrhZpKg881e6D9DbuRIRJ55Rcx
5A99VrxRbNueX0QVZFEFw7BP8NAB9wC4pHf6UKTzbfPxm8+5os5SJGILHkjBM2BvNBkeVuk2Ok0Y
xKXhqIc5zyXxuqxYoJt+SkuOeCbE0YcBZEP9JTatIEjizuWN6nGtYsQlHDD1qZ+/YOM4zZOYQN+e
PGc3x1P9WSyZj72bV067cp9ZeFa10BzfC0SqWE5+i4pBegn+yG1BUgs26WJmOoOWVoXrabf6/EKB
wzaatVqkScosoNvOIsRQG1N7xf4Pt5aJOENiiwyZcCI4jEzNDha8sSrIStpFeQmp0pXPyhUT/tq5
q/4WdN0JhXCmqfvno1V2awVRBxKRUKu11DFuExxOjRR+8YDls1lHI2eXH9SVLErxhaNxS/XXZR4n
RHoVlvEByIifqFTiYlQqwxkKehWAvLEuKzfT/L24YG2nRzgjAzCG3pNlACvEhmCDShSipte7WW2Y
NCM6HnN11zufazi7ibmRnmw87YVCcvSy7Gyvmtr4/pH/4qdiPjg0MDoc7oJD7aLoQ5geVhgqdIsC
2DhJIwL9T6HBT9ovzkzK39rpA+O8U00lQLiJaTmb47mfrQvt6Zaoy/x8VXl2wA5Qqm5H7EAk6vgW
bVpEZlQiJ8V1nhnUYJrH1RHiaqNbGJzbOpI5MSegaxR8uJCbXDNRvgEPYjM8qCfFxF+3SiYfkAX9
EFaqiAd2CQscw4G68OoMrPmeVanu9HqhsPcMcDMlcKIekFcuTK5Cyo38V3+2QMdkIqBsk8mfbFqv
TiJZBtcIXhVhFT2L4GvNHS1exIjrPe5GaHTCYE7OtXP5MGuqAQC19h/RgpljC1rVCjOksKwfEv3f
Xu30Z4sWiPZNhr3Sr3FELuOhApHIGzC1aF4vRraw/j9JSUFFuG1GvMdS/3pXT+uJaM3rH1FEk7BE
Ru1XlWJU1M1CXjux0yMP15KJAYFkPs8s4BZmbs5TVeSRv9tBTBcKF3gBFeXnclK5bPXqKmspUSRo
xPeE9haD4Tl9+EEJOym64j7C8EX0hZQCZ6S8TobMCeluneuSeYjQ3cu7uHv/xag73KBssufEjM4G
K5cYB6Kb57JN0PxVqK3gtbuZVFCWpua6Kaq+t8OOm5djC0WcOC2QictUHqKdPFGh5lI8vtSVKQyZ
u8E1AiREu6kWpg64mAK/La87ZCpUR0p4W/WRbh6UlDFfC41CchkSU/NDU109NV7Vs1HIHfc4C0uj
XRsuKw0qkJQ5XiYiURkjRSptLr04jTDkqiwUnMAU1+12AU1QCgkgKOpV16JDzYx5w2MGda6mlUlh
bBmrhsZGdon+DYpoQoYJOLHC8Vq+W7lZBdfIi2rmtH24hYbojz8BuFliZZlwNzqe0YzAHjm7YUVt
/VNYuMStVmqs8E6C8MMNcZpaTPpyNimmRchV6kosKrwUWtwYkFKNnbxbG3P8UWxC8FzP9kxvPLRM
HIxdQgBPmxJC5/HL41K/BWSF9MlOZrenbQpv157GA0IqY/rDuB7R2zSvBrNWRT/3epg91h1fs0m5
MV5Y/BSWvhhOfzAy4EDLxe3tMKjXhWeOSd5oYKIlDsmmvfbTxQi3mVOTmO/S5VCfFsjlVz0hNL13
ed2FFFaLFLgVqHZDBjCLydo9LwmXAPUrzjA7Z3e1tx54k5ngeHbNo04AN+/Tl4hfRV2nBTbWRvXy
vu1sTSte1VAfo9EpymWBEHgdcuibQyFNUs8wwL632M788dpQA76B46+I84iFVyY4ZQXHchgtKqr0
1+FjiBfVDuCOrzD/WoAv4HpbkIfldZCh6XEbIO6cpioWSPDTPYILClq1WpOujNekp1kPz3hCf7Ak
GsVcHS2OWco/8TsaUQCPK4UhYygWHSoFxueQxhwG4dowLPNTiyRlGrCn7LHJ/bxOgQQO5RXOBAwC
rcSeipHGCTNpHRTq+5bw+Har+4zC1j4JPVHkbiAYO5Z9p30nZxIo37/BY23El8g/K4bYGdARb8Tr
WqZQ0roNAtxbybYRiT/c2ZGFmnA+W/ehSLWs58S+Ie0G7KeS8WCwfvwcWsOggrGd8A4YOmlp97cq
WiXKpN1dEbHm/XqPIyoJoWfskh1t5iKEnKc9AjMGAWg888MbuTbCHXGOs/eER1LPkB802C20pqOy
icsUJw/ZEkJyGpdMXP3Lpg1w8yur7zLpJfQJ/YV1MPpIg2tYECWn1c7FBhJv/rc/SRQ0770wez77
r5JBWmWXkh6haUO9nqgMc9wFLFXPCytXSPjXnz+aJqViCD/ZQQWI2edVx04LH1lDXP5cKZTVXDba
LYbjg76eFwiCKPgytendNlM4OPy4YQSiE+VC+OBK0pjE1wZ9WmdiGnBUY6DQ2hto4hCWmU+L//yQ
MC1o2mF3YY3jl4mR3287CN4Og6/S9ZqEpAuiSlrMWZr/SOXBgZjzjgNBRpUMVEs8Ell2hs91WUe1
uiNMN5PkGKSnH2zyziIO5yV1VsQTcu7HHa3lR4zR+myJH5TOk0hqsvhwVzeg9MZV7OrBb2CxSwuD
u6qogsYIuWJCEsTdmEyYxtfE8hKNvQH2V2lMAGxSSU6JqTUJCMkqLqqAnSwUkvfIY/Oy6DyoJ8Ue
UtiicRdMWpMQ4fCtQ69cWueRCOL0B/OCSqWGRgCOrXcfyOWvifFoQK9IDpCK57MHaPlcrp70FZYk
5pmCupGt/1IYBbkbe+elBCsw39d67OSH2RQtfByioopc2nl6NSyebvz2p5kCu1SbF6y5rpaRf9sW
h3WfJFLIW8ha1rVw2YXaTpeyN7WEPphpu7+/97BQYMw+F9aLMiHs5Bw2/WSLRLpdgsbnBC/cSK3i
dpxdBfcCIvrESk4YJX7m1pMD3CI+XnS672vmooqv2TrzHAZpx5LjdbkMo1GJKRtQx6qfFXWspvxy
BqK4Kq0j2qHMEvDU60LmMNKSvrjfSDBe/Mf5a/FKHOtTuk+1Rt1x7NG3rx9PwViM09mUDFWerYBY
/vHc9ncwEaW7aA+I89dA5EawV+7yoPXToKzXH9iYLHPuya4hI08eil8ghc5HII3m0f/IcrhIRcG5
eyZMq/bEbFRt73YaDSucRyG/Y2Q+cyFMgexPiBfN4C2DvcyAmaJ4XITI4Rsat0HyRC02RLeBTMWz
6jZ2lmLTMJXqwqWQQn0maHSAWX0qEWUMCjsTGlWTMxpr3sufsoSM1VnTW3zr1GhQgbVguj4IV2nj
QrltCtpRYR9J4A2Hti/yhLvE0FWE/FB7nr/B9wka7TTUDUBeCP776Z3pV1GABoWvK8jGqKUprdjL
nlekwQ6wgCBjYK1jd4MqkL96f8imbK4sCwqaxwNXCUi/00pKPATd4J5fqS9WLLiCUxbX/WAwJu5H
ZAEmfitHrxD+Kif6WCgBee+cmUwQoOGsLbp+HsUprld0vijWcwN3zx+iuXO3IOn1k4rPnryoOHLM
obHltewpbDKtFB+vDJVEkzFZxaGtIkwOpnX48iPIWZzNGqyo4qElvoEKbNtfNQhj2Oz5jHKgRTni
AyCxpXAhyFRves0yc0JRu3Q6zjM3iOI5J8Wa/t1fLt2Yv9WTbTKFIIVMt/xtigo3gUmeV+lhEKHw
9XAhNwINPr70vqtqd+HSzzxN7b8oBTi3FM9t2zCfPwkp3e3XRc/AqoDU5cX98QSt+zua/BJZgWfx
G1gFpEhFRlIYRP5SDj4TYuVXwqg9ndHO5hKsl8yVfCfp0LoyGF9LZBK7Tw+vpBzeCEDRNYYU4IAY
wyJ2tt2wm1H4CDcEJLwqCfRnLe3qsNYxEDOOqyZflMXk4IYKXlezLoi3vpx2dtki7bIKtUzCR04I
GxXyB3TcIe2tDOEGahj48ApjCcdJIFStv5cXRGlJkUEfkYDWdPcXcWluVu5ILUr21iVcj7Z4dwSY
Gkwni5RnyxhX3iyEugJKFo8RkuED8fRTNZfN6LoLdowT+izWZ68OLwkKCkXTad8R3vNQTmkn58uj
jQLniy/1fuOKsp3MXqUtrnkYxYuyZUcYNmyKLLY8r7YEXj/9gAUVmtAdz7Qi5YuNSpQlYYWJZw20
m3RI1QpCf1nUrhiqBVU95QwCvbdbzAasOfgDQUMBLTPVg2o8yxtUG6vtZbiW4UDSISSPFMJLtNiB
VB+gLgyskKWRiPtNGgwJWkn2A/38x9+4YeQE9bctddDuHlk5mH6bOxDoXKUAZyK7UuAw1FyndiKW
znliRjDW0e0G/WplauqLI84QMq3+EkwKrOtVCCIirJ9HumLWLkk+H8eTafQ2CK7ODlnNBo2ut0d+
+W6w1QGbRxYIfCpufdCSd/2AxP/ygN3QSgTJ1qha0kMAAmAyQ9VNeVzuFaQm8EI3mwFdiDAKYtVd
SGFSeYkggCwpzTeqWSQ9cnaMjRypH8F9p7WPt8El/QpehmfhPAhsxbMG1qIm2J2hOisV+yRqKNmx
GzEZcSMC5/fIRlB2vh7O9AH93OdVuxC/wfTyvme2x9w6p5/Nbnghmad45i89ICqTIUjvbUS9utWW
QNa3wkkBSZw4oK5HRDLiqS09gICdzEfbVg9cK4Rg4kg+XzgSpt7FzXtR3Ilr/Lr0wAC7Qam+QtRJ
Lw9eY+MqeI0i5JnAO/XLb7Jh3nylX6Den4F0NMlfUcxzvJVzyvWAb+VkvBvZZgE7bJIdX3eUNGXx
FgT51YsPrj2IwTn1zM0Qoik0e/iuaoM0bFl70pj1pJIfd7f4zchkKUMeNGPAPPLr6QwvvmIc7Znt
xDHp7UxsRSvac4SkUVpzA21ZWNAr5ylNRHQdYSudF/F5jiaOkpN1AZoslhVMijfOJGcqSyVzP+lV
PLXTrtjFxXfnUY31bi4J8dqqwRl5ydu4CXgOW26cAzxi54PR6I4lKeBOJAlvIdXS9CSgv6GoKQhj
zfo32/vC5RYbeWe4fAGim6F6k20IGmcag5cScLVvKPXDWZEu9YFDw4KWKi0/+vYkirQql2mST1iC
6b0A/Cj6wwbgnnSuC7JEjTXW17bvfk1/FMpHhIR+JHmL17wew0QLen41IZOlMWwwo+8gAxkCwGD/
9UMBBL0TflCZf3vcKEGP9treN39frCjmZDHFf06QLcuL4Oi3R49ABrx/d+EdqLsJlQDc5Ca5Uv2e
c+GHZ8bEXaGFas78ZSunXI98JB0xaHEGe5Fdo7CBh6PQCEeR3gTOOJyCLFeSlg8ev26s6Gdg2roY
EbC9BUs2oSsERgZ6tsEij41vNlSCQO68++O2uj7KIoM8DgkwDmndiCKXWGO+EHIGISmYVKDyDT2W
2eeln0NhS4k1zwqD0r4F+sACZGpmzplWVhLujoEJgSWDD+snjiKVnC6fPNsSYlwlWgzWTZIMXwrY
HsRkkP+L1+OTDj5B95EWJTBf/PeVxxBFhD3RMWNw3GqTqJQ23VPJpSv9/LGCxd8UEzjh6fAxrcmY
VqYPXLVYg6SLbTe/lB7rI2t5Q3P1ZCWMMh9DOVj1uT4QYD/VKtBS4mRwN2Hc9VvUnGowTFNY5NPs
Z5/R0eSHnub+Hy+d7qpZW5r5lHTcNr9Th3YNybowxJc928HyGWy9P1p7TOCZB4b1eqyVUmNkFBd5
UWlq8Unyowv4MOesB3mXnkvI2PFKm3s3HMDLlhrN5BDYW6DWS/ARXZDed7CFpnMidQYsQkk/yDpQ
d48CvjedSImOjTYja++Xz4aaTyGTkNojOTvv/uX0aS906qyGyt+ngo8724QHR0KOXcjcsfelmRaj
PjDYW5J7wmG3eCO0wiPh9VKMQSTRNeQFQAQ+glEijg5XssSDAYXJFefUGf4uCE2UAtCrYQDoPJn7
nk0pL+sPu07udklQK9nUD/d/IMxf3c5CVJjrn0Ut7N8GKdsDH33DUUADbtzbICAVoRBcz6vRCLv5
+Nlj5UcZAfuYrp2/yxXfKUXZIGpsgj1swwgoaqI5sO5mDCpCcSnSoKKXUB0c/jPISzsDKqS2Ro6V
rnpzFOUyK/GAr5/7SYRkJnirrrdPo/scmeInSCG8g6f/CCDc8HN1tMf+YJT1SaCsaCecQG7FEgfm
l28Sod+3YL8cASsha/67xdkjRo3WfyFIdOJM+QV7s2WCs0fkBF6t6LpJRmdtkeQYq+3qPu4yexuB
MKv7sn4jRetLwRs2f19d1vJndTR5LkFPov/Du96/W50KXCTzK09QpbUr6MIXuqLAvl+FguRZ6u04
hvOiiW5ydSskPUiFS/vk+EXKO09Dr7F/z5pNfKycqHvi24kpddQo9r5iQyrBaJHIarPgKz/Bua9M
q7VK5hbQ7M6OqwkexNjxIXZ8G9nV//wfOZURo8ljDeZun2SipA+IMlO6U13EVaTEsOrJAJnkhbQR
q7yZnkKHWTIC1b5j8KrTf5lg5qdNMS/e8SAhsUeTHhl8bpSj5A6ur3zwF7c9N1550aNqZs287gm9
foa0uh9kX4uMytoGY2CNFZkZgOaBjrhg64ULXaiFIj8Fjn3aN1kL/6z45Wa1Gwlg9UjJG5wR7KE0
K0ieodkXItlILvMbWsuSTlgOqjY9cwx52W1rSsztl1gq+YWCIzz5xqPcr1CK7Bz8mF+wjncUQ82H
kS6A838X7CsfO6P5EAOE5GQQ7TSYXXgGfGgshsDrsCGAlNwVeGIGu6Ur+GFO1L4bA+69lbelVOsT
uGmaVoX54wDb/4hIRZAZVgFq+tpj7TpGUx3sN7rHtFMxqbC4J//B8fJnFd+sia4hiTTXTmmVtUfE
YMpjroNhJtfpthuqV+UVVVNkfjLnSqAyTnrJaWYo0VxcDyNXULUB7kdqfqk6rUjFSIiZvzsHA41P
/vl1D1RDsTnDvPPVjponqlqZbY7U+ZWHfrE7quGBUy8vsf+sTRcNzsbsDIQAoTPDuOj426erthc7
sc4YubGZWr8pp0uH6Ay54gugjaWBHMWD4dZbHreDt6r7hhsNFKwcR2uKKRZYO9cvqiMdtSW1h+YF
KdCskXrgkh5le627SOMEP/zRwE3kfzqXbP8qD7qaUxNqZCq81L0MIpc+WDm5q44cbbTqnVSNcX9L
74sHT6110y7aVQxu3g70WSP1IRkZVGBbMdIqhgyS0x/PAwkuTk/keqOJ7QvTiJnxpbhfyijcRkBi
dmPt4PyfrqObJCJbC3bRYog6c4DjgyAENJCSdAydlN8N+b6FWlu8zT1qSmAvS6dVRpSqn+f3PGnP
zeHWnMfScU6KR1W8rL0GPIWhBUAqzKPX4EFZaCli3ly2q5kX5Aw1mtGY5NSmIh1mgRNBi3UKi++6
UB0G/4DXvdWjA+X2AKfO/i4g+jH9lTwdNCC9mYgVSu2UXJncNfPrgsWRQxfcirwd6PmVWoBovXel
BksVYlQLmja4WPZUaiDpZk+Vw0eQKHBEd3s4LSTPailuN/O2poe6cECr1BRT+R7cdTd0SSxhsUKa
WWeEvD3X+4oAb1RVQ9VNp+a2c2n49s6KSMf8tA6UHLUxqZe2Yty3bo/23k/VBo4MQeV1YwXmQ9dh
nUViT1bYT+lYho8Z3nVFvfWvPwwJQtOZ3DFi7KzICd/bvhXP2psWkIcZc/FqY3m7UESXuyBJtLX5
b/0W7IVWaZ2BQgXGgo2UMGIF33ZVw8pUziE/r6eBvllGbXno0t7gKlh39T/2mGf3BD3SEf7RVNFD
A2jEw2nyZ+eo5wy0DGujXQI5xRy9J4RnZi4WMNLltcflYGcgmSUJcnmxALE2Q+BgMDQwstbqDnXo
lSMylkOmBjMThAi/82uPVrucd2aAuoNkXAVOzWL5tEMXCe5BPr4pYyv/XdCV8VmPkAvMcHOC+ukR
TqieruwiEpatueYe+sL0y2oClv7/XEHYmUDIQDVZ2sfPFz5XJPcGnGj6j43KzW9es3xnwW037Y3Y
n4/REOzc/9tkDpsRonmzyzalejuW9vwiyOkzkdEOOcieZ4DwaIBGJdYAWDZSuzpsoKeWNwGvfbtQ
jhQfQkRw199sHX4GDpCi6kImyKFOsq/6eMP1SP7Hm1OakWtPejRRylAso5gOYh47+DLbxXBTqXcE
mwSTwDQ4vBOn00hEiKfn+chGLxoOxT23gzj1fm1Z/6DrZCY4Esz8xKNvWIS/f/ATObAcoP7kUCf9
ByKb0EVSlBWJJHUOaWp9jHVAK8E8UonW+BRVQV/964ZFvJ2R/fpQL9hrJU7Q78TQoZKKLi/MLwri
UvOx9vrdmeY7qMIbSEuCCXhT+kC3FTBLn0ztrzice79F31JeUMu4hXARLDCf+EVjpzn4/VIjwg9b
4F9HJPK1oIBqvql+dEbRQ0Rm6FJ19ZepOOVxhi+q4PSCHkpt1CGuyYiQi/XSX7uIsyur7H3ZAbRw
AppzNtMxIQ6R9N1DhCuAbazwOK028ekXcE28XfqzulX3RACbfbz4bs9FlryIkStr5sEGl+8fMHTu
+UWWQ553S1TaLwylmhC7rkEL0Zk2Z1TsYH3eWOEB2cQ3ez6yg3JD6TaKw7IFGDQJq0pi2b7OpBsp
YnxKUBsXxvLElerHf0P5WgaqfB080cp22QX5W+hLdXmeN6bi/WOLMaQKGhr7zAp8oftlpnFH7X/v
aV7V4Z17weOo4U5k026sI5F7ovmyHG7BSALnWpXRfCmewUxtkhDxEsx8D0xXIBfqvukHxQhGVG83
TNnLJCvtyCnHfmmosvBrIdJE/hxCRafmuamypMBEak55gCygPzNDF0YWgZ09w9B1/PCXwPHRqqWG
vKuF+6PSkJ2gi7AMoobZ1kH+c4svzBfyQGMeECaLeK+0vGg1oN/SrUH1X0HaGF1VH5FUOeWRwJWq
0FheBeTjzFs9MEQlWbdA6cA+m6C9LzmvjVpQGIR4J4DUpUm/PzhMufy0sXtLs6L6RStUjPThNqLL
9c6I9e2jQGWLAOOhRoU8BH9ZbwHqJ0tLUDetGVkaNmUpQfW8sKtxO2qBcA7PmqZ5+B6fnt2ug1Dr
d26yit28Yt7tMuNNHhUyLrMQ0sWk0Gws/ZIFelDt7Z34bb64HpXDUXYZ8rHzutU6UXStGlGtgfqD
gh31/xJuowCcCXB3TIO2LmHlJ1OGBiNXaMbPhUDjbFVQkABmxX98bMshYR4KS7Fb94P1W3LP5UyM
VKNG9GKWK4vPSgn0soSRcQCOYV7t9qDKZEi8NslrocJvMkdVqpYq8v3XUcjrzwK49+froJ+k89dc
kTjXB+6+Ty0/u8z6w2TwPWA1CY2u+PkEzWNiQAr24wbU3rIVxZoMbqHt8NXzSAsyo/jnG4voxO1E
SbvcyO02WMxq/EMPGzTVdTGQalkTe6OK/fghDnWkWu7i8BiCF49shVImqJ2fYhczTrXE27qHYngn
IsLRQ6RER9aWzcM1SakDbA+do7PZaHyixCVHMCnE3bruDnONkTozpCQEjuJAGqVxyMBpjeuI16UC
ubkME7rFhgM27D9pWc8vdumbxkM0fLo0HZ9ryCDFGsEylAiYjDtQwLSrfuNOtyOk8ddFOj8KbnE2
70SzOnlxw/kyHfI5mOtF5Gvttm7lbNqT0FwWhlpvSybEzzmvruP3Sc4AeFgBNgRS3VFcxiPpChes
8SKUv4XMrfrXOyawH5WLS7CLWQEt865yyMIoAMTHpdXphSCAl6N9gOQpKa9rIaJNPwpzD2/kh+en
m5fMMdMFNnirSaLGQRm4M9QVwZL99+3moYGbRQRSr3oNjIDYftAg6chRhKKB/Nq5tJLRjDpHsrf0
C7vvm7ZnsRTBuow3lhiYm5umTokADmi6jIKPNj+uZ0XmMYLZnqWBSusWuSELVxSPgLGtdmecGIpd
ieDuJuQeoAd199r8SrcG/W6XlKY7ztAE9rsl3wKI5VFV2oKOQkQptQZkGxAnuawltVXxqd+2i4Mv
EX7RN+VEuNL4USFx+WgehN1ZDtmIf5NdIrKuhnhL/SHwr9jh2hoporzfP4Ol1M26zS26whSBxKga
FFb9xK0jDf452Rj+r3Cw3NVS6Bxv0zyteajvSSJkw/5Sbk/kGg6b3NLrAZWp5XUb0XU+gQprYlTG
DV2zBot5uOMP9zCeyS3Bw3DeGYGtqOmQ50e+ihWhPdb48+VvFci9YTYHfkRgdQNnKAWJeKuFSb69
6hYfpfutOiLoCGpMhizj2rJQJR3TiIW/Fc7rA52VPVeb/pErF08JGowzAdqilm8ven/ec+3ug6/U
c093gDZSS0IYUgtjR0LSW57/0i4FzSDdt1ylYh+MrCWfQ7oC+fFqpXdybGxETqxR1ZU5h+ie2V1Z
egd+aMZeyx/b1X+LI7McJ+gG62IqQbAuuktVuOJCTVefiEFv8DuDWsYIESyvhpI4hcLiVzhvMcbJ
SZL6mOEzBxy6rh3McyehhSIVNhfgfFUoQwB+YYmFULkqX03sK4y/P4tGMk5CCiVFIWRDr4NHIN5h
mYL3hMjBCJxGTw1x14k49IjhunE+X1iVjJU20IbKf1/SwpSnghWfcCJ2lVHwBvhzbsP4/3uuU5pm
2IeQByaaSrsv4jQcuFFH5BYh9LWiJbrBujwcZTfKF8Ly+3OTgpa6cRtq3X19Y/H4p7MFPRE80Tg3
/xZqRUUyKdlFlmuL/Rh9TcYTmtPRl4MBVLJANKp9QqS6n32ApM+oLvbW4PyO3FLLEmWpuvYFiSfA
NfknN4pcXvXRDcaIh3FM3ZqmvIvbQm1IlMtA9SMD36dnYxdASM8R6I4Nk9u5ZdbpkgHJsNu/wk21
WlVFOZPUrJ5UsSix1xHTTmBSPkuF9fEyNG/dCXvMSYuHdU8z+eZK5rjivFrxNsos2bI+RDHzYVsl
+VnOMyZjc6untfViK2ZN9bW3D3Rqmp/1pcVtJPYgNiWF7xOX0oi5unDzblUoVjulpWgKQnT/dsqj
tk6GIVNN6vNFwutWOoAc1SEnkJnalYgBH/HBPqwrJPEjvYCjTBiLgTEtt4l9Xf4dz8mU/wQqybd4
hRKl4arMo6ni3PF4cAHSK4mgpM7oTlONexRiEPcBFPr9fREElKrOMJH4M+XAqFjrlDx7+CH4Oi24
LPSlj3yDr97SgEwsYz+GqzizUizStRmQFMECw7ZiqEzcuglDoPch+VTRQtDPY8Iml7kYLsasDNsw
TsodAGzwK3JmtcjJuC0Cf4w1g8tIVljfKSffOv0kxhDknRrM9AUtmsbVI1WCF1zYAk08lScZw3z6
tQctz3ehpp/Hxw44uFwoibwsSDPdPTNQSSw8d4r+blNT/K+hTuDtsO00125wqyhGJKKmHQ7bgn0A
c1/L0tD+v5qP0O8VcW5+UN6ATi20dyJpsS+4yaLulUicmgggTz/2VUb3kbyR95GuB2wCwBHGNI9j
kfI43cFaOxadjTspQrlOCgVCiFVGQDxdPonHA3OYKkxYb0rmxqiPwJbC/Xkp8C7fS6YQykE8I5ha
AeYdOGTh3MOLEQtK+5uyvThmunhpoYd9G3ZCpP/Dey2ePvuWGinzn9d1EDHLd/lN8HzO0Z/ih4XU
nUepRnGMDQ+2XrpFMVJ26EkLCPq4BTajBS3IQxjk4eJKkh/IScdsEsUElPDDo59NM3VeGrmBZ4Um
kpkuFlb/b/Ly9Tt0Aj1FXCkovfp2A8CweGZPcHbGt9Z/E+wN4fSa+SY4UM3KGXqJpI1v8sLaj5dK
P58gY7piPtcSJf2pShbkxPK3V9pygWkEAdsq2w297HSB9vf/vKz08mJyAyQD06MY7zXSfoVi1fFF
Yuj/+NyNXoh7qt0R/gBb9oKArnLYSe+hTNs2CFFUmIggyTW9+S0Rg/lVZtqmlQbHIehjmc80ITe8
70x3D/AZMJLcvAuO33srlSHs8/jMne1PUFSWfN9dWSoaEiySYgdIX3HhJZkW1YfC4Yea80n8gGFa
BIUI5m2NVJ9FrIbmUM4cTdOlH9Fe/Yb3wkR6Cq6tGpMs5geh9ZjFs52eJv1pmnziQcs8SIYChrRK
x1tG5ZEzpxmyS4yRyFL5ny7t+Pyw8JP3kp5jlAEt+M5+1WiHBWTvaHP6uCJX7g33349k6OiTmSdY
KCNgU7ypDsh2e2CRXUvZ9CnHXsGR4gur8aGNZ7hbKaNioRWh6LcrNkwTdESa0BGw8fyEFhRea+Wi
h5RusWZ+7Zhkaqr90dtVSvv55ezVs/27+273G/wPLBPXeLZBXrjOEAkDY97ywuhcNtuLZsO8hKqn
2Iqnh2CDi/Gu61zr9ZvTpR4rzcAkidZNumOSgZwWMn0Q/2780eHJSA0puX3YIp6C5O3NEvZSrD3e
E8nIq4bUdejoG6QIdjoT+HPpELEN0e1c1oc+SJ4Nu/MckB0CEes39TNTGHaag0r7615tfURYUUzu
/3HPJBOSbLIBLu1DpmqLsyLjAQAlCQapJIH9wCzmWoVK2iNnQeS1XFkhinMWeiijWAEBZ5f7lfAJ
/BsNNaoDWAWnS3SZz2iYAIW16RtlD9RyaJBP/gJLxkOnJDAHzwef56lX8XojhT3Hg4K/KrFndQP2
p/QyZKR7J+dB1BAr1M43K8Z02TXitQecR4V6xADX9Yooo+ou/8SL2Y2gX5cm90GYiGwgTr7khTin
eegRzwZWr12sTevU4YnBPjCxfip9qX1c6W3myQggYljPHHBz8IEG8ZcgDilk/U+7nj60rp3AyO82
Ot9QGmhPxS7naTvIa+cYyaMDM5Ft6SY9tuwUOF0Mgk/+rOwcq3/mP8nyh6G829D6kBkh7VFtW1ui
EJM3BOrZC4mO4WwsQKwMmRM+JO8vsSNH0sOUKyyUYeG51YBnI43s9NtORd8fxlmGNEvxk30i/nFh
T5is3FLansU0UDF2UvnXysX0X0BMfxbH2FwhJSmSq03mzObqqh+4/wwAAlfFBtfHn4N+TdKQJhtx
UcvwIFl48WgRQal05IdY8D7HxpmAS8R6Zee7xJ9ICWCvlFM4da01M0GegHKGyWPTNSEBRKYnBlQL
3YIlLVHXG5A740uE++Q9r3gVMmprvZ9pm9yKGtAfRDeCMXc0+DoQ4Pkvodcy7Qj59ehkTI0KXd+k
EjpwSOUWOXybxmIv6A9EHBx3ONtVmfOyU7hRtJcOR3JtXQ3J1oeXzKNSr7mPIB8NXTQ6G9mnoLr1
H6vVDrdTGKz3SD872dpjF0bRyypLt7nxJ+IpTTXo3aSR3+xkz/Du8AJfGpE1pBhutf7tdL3gBhpH
9CRYoPiXyterTiP/pdgFk8vfUFHG2kAE7bbuHgand+kHDPqX6Cpz5WLz2fgMbX+oEY0jE+8+kbej
hN3g6fEscpv8gvaNBxybjb/ABhX6XM1WxyF2QXpg2SJPswpHNm16rCpfyijRH7fB+2woYzSINaj2
ynQBFvDPvEPb7foRfKhs9g7LpeLaJtbT0Bc4mIr4qz96SrPk7NVgqfUz1eX5fGYnXFFPXWKwxEhg
K2VQ38nME4SybCLufII3OowqKGozsPxOLZDAwz83PqqLJtuve2ky6PRgbD9HF+XEK+l1SDuSQGTZ
uPHP28mzNCZ2SRS7SWpEyg/dReZSPGlubQ+QdeyH85j3sA8qqTaPpAb3AOoi5cIe55l59q4hbCrZ
wjHIyxIgIdpfSYWu/eXxMuN8SYSL5/nTIJoEwbrf1l367iEB8cecd2Ze3OrvYzIuSt/qmi47ITZO
MOnW/bE9zpGA5GnzN8RvDZpjYjoG+Q07PDKCn2oiv1i9TURSU9wPhUz/m8YX+qpwT3PSY2cm3U7c
FpdNAhocTG/x4IjS61kjSo+YMup+9kuXqd0gBPqfKR0pJTXWvoJ5FZM0j8RRy9EvtFZ8jWrJ87x+
LGY9KE285AKZnDzh5B6llr+ok763kY75RWRKwyNNHGWJys9fo+7ausT6G1AjdyAPz/0LsSvbQjIM
HORQVpKT7gL95GIOMvHzcRv2LrUzRWN/t0KB6E3yY/vWVeYAj3HT38RqU4jPeF7tzLApQlINI3wW
mp0RFx15nnmdHCLE0ELUgbqoCNFDBUMTElOGVShjjHJi81VZhbhzxGWwc2X0qzyPtX6Lahw9+L01
PjXnBhX58U6pKeCczb4Y5vn1Z/uU8N5rtKpW/zrmLPrrnL9df1r/P53obJ8Lt7g+iLYtMpdQwVnV
CS94iFBVMNhPZ2Op/bbp9wHIRXaMWw1PFaEgISXzs3USnD46VLyme0n1Ph4i0OiitxXgrk6nf1Wn
P3RmMruv6jB3h5GzBDTW6/jq9qAZ7A9ybqaCvc713D/LMhmocIimeDT+5Mthj52oK2FDb6uN9Xl4
sk63QFwJIvbGQaFJNfuf7wtNT3EpQxnGGxN8bDITN8jKcNnDGZ4qjpCJUewGY8rWDIUV0j0IjyVK
zhu76GneKFu11jqddg8msw3lzEgIEVHsiKNc4AQ9wguleWhobcVScx1xJ5XANX9nEgmRYvWQxGSO
cU/Ut+8KVBlgwyU2lD1LmL920eXmecG4WqAoiT8bM3R/3+4tHEt3iSARqHQ4lvmCBVQnoy+RkFNs
73PXfaUoBMiXVMcF2ZP6SRjTl9SK4ujMLmIGc0/6L8uqXQq5jAvSVLKIRQOzGZp66M86/lfAwmcK
fkpY6zyjLUuZxKq9O6qwMS6bge0naMZNFQs4BKfdoMVexqMBnyueEAdfJTS113ny5uVmMGbAILj6
wEQVqhsEikvwzdxFB880Mqhj8zf0Nc7SolP9/EhKkv2uEZH5Li5xFsXnHrHWyjP9WcxUAB6cYaV7
ysKKl6M+7pnfOksphSDac2NdtuttlfFua2CR5qpmNJiM0wLcXj5nPZhiOkbH8sg1iJA3uJeUwwEj
CyQKSnfpP2IXI90vmdwO5ZM6gT6bkgU3VFDQHRO+1OaVIp+tKXO2hhgSE/SNjEZaFCBCX37BCHI/
JxP5SlTlPoHXZzGCneorUewq9abYIXD7b3mIj5riz4T5sgQITTAyQT6rfA+Fr1xmTuEejAzSpUcl
ZQfXomgpBwGUKCx4zqw7321K45TmCBbYfxLfCMfhEAvyoXUZBQZHU9f36ch6IU/7Aju9kJKHv8F+
m1OvVErgJPUgSZ2wF23F0yJwjNjMCPjQ0zi8oTJ+ngXgkq3bdPxdcNNLk/rUDkNO9kHxudm7TCGq
Ql64zvRP4gD1vcPbF2crMASlfGUkciIZfU8Lqsq6vcvldCuBr4zAkUijGbXdBeY6f8ng8vgdVxba
IJ5Q2wxCSFrc4X8kDkq1A2LuRv/y1SQAUmf6J5IXJyIZq6x5KvjunWsXeCw2Rpz3mdzk2LA/UdwK
Xz167+BauNL+ECyb5tvJ9nh/Ksh39IlzlWg9HQxkTKn/hec1lAC78EMaIlaUwYvdtzS72ZYxfjBZ
6Yb6CtYg3pK4lngRDTYKW2+3cjnmi6PC1oW8gqpInp2OqxdF4QmSucp3DzVEFOaF6OOgl37AJ9F+
FJUAT1rKQpVGGDMIbsfgJtw6vJzl4QDzhQ96jSPsD61RRO5D+UtCy6Fuo/8noCffU9VurI85quyQ
i4MlxOfgu0iggHwQglqGs7GSKjJGTSTEUK5U04OgcpNUPli49/r6edgBcr14iQ8TnMoy4H8qLAKX
HAzYWd0hWSpRDoU23I+8MmzKeb5TbdCb7Ncq7qCCVKkYO9xU2G8JYKJPZjLlVrwn6SWDnqY5/Lwg
uFOjMIQSzNDDjSfK/dtbg+G84e5YISO1Z9YSKxsrModsKOZKqHpQnwbpCPv5P08gcneeGQ/qo/1X
zaqzw+eSFtIqY67Hw06u2ScZvPa7ogD4KeoHBmbL54xgDtvIKAGDGAM20o9XYUB3LDNKa07ngQoV
sr42MisGBB4aPc1KX05pXo6mXfggUaV3aQeTMZTZQaun3VkdKbMl5lQYDe9eNqIz8KW++t2fPoNn
9L6Q8MUuMbX8iN4WwPJiiCoC+zvQxGt+bu0/s5XPkD/2D+C2WEe0xWkezqoyrq7/jiklEFayhru0
pQyEN1pwe6Af4JextfGY/er1YCAg2xDQdkdeSYF6M37w0K6N7avfIAs+TTTrF3CjRoaLq5lVGUB4
ywt2ehnTIbWnbfB1zbDcT8qgiYsM/fCyJqgABmswUOING4gsJ0cK++0m+SLTK5IE+To/zgUwnq1q
23k+oS5m+3zn86SCJqGZHB7NToWM5nNcm65jngYTLQCGIi8C6wCsPt3IfQ5BmF8588cgZh+dQbj+
sjLix+xL4BwzOUPf5Kx3clt3WMYY26Sr0GYZw2RflsvNeDrblWoZtZsVvJvXWQUSsbovQ3ToT54f
9BGB3s+uLIWWexd73Nab0O666nv6KvevQ1SM3xKPoqbuXusuruN837Mo5/sl4XjoXVZSNPZQxREb
8D2MfDH+mIKupGrjOyQM7UsTe/i+jBAjh+RMMQFz1JIVcpGZuQMJn/1hfDVWJrQNlz/q2dxY4EL1
zVNKRtc/Qrp5uvwn8Yfa3FO0wtwhN96hOcReTHZE7e1ee2RMp0NWcvt9hxv0ItY3Xd0fk/R5P66c
KLlQojE4VJBB/xn/4Zp6k1A+PDLvf5mZFphfkl8zMAv0+J97Zcm/bSQ623I0MKYD3RtTV3i5Ovy1
Sb7rryhOK4mqg3NPMeQWN4vZiC0zCsGZ6fIT+VQNj44mt11Xc1Y2mA97zwTeqd+hzI3Pgm6PPfdG
DzMS+EcGmTniGwy+8sNUnRcRdfpv7PSvXH+r1fTWdVXdh3CylSm0HPNno8A7pSyrkBSX5fxBVKjR
w2oIJR+a3WucbRb7nX2XmSlEFt53khgJQoX2olYZOw3zUFVME4PeH3xeXUmoHIdLP44CRz1DQJZy
KUpFoD+LXRyJTMpqljnCcquiKfFAN4B+B9RRo3Eiu2ZWKYg0GI0E3NshCafVrsbPFkYs+Lwi0gar
maJMXIkXcUubj5IjQJCoDDKDjzHKnH3NMP8CDKG6vw1L9szqf+ZYok6tq4r8rBmq5hxIPVlyn81Q
2nOsy4BIt+pmLii+1nLFmh4kWLqpDJpVw0GR49c0o0bDEtqbSnwuXXlAiZHWtyLqc6PtHUh5ewMS
hCbYZrxvsx76YokaJuNFZn0hIfsIliZaJjXAUGuVfFwMS14pggrtDsDokYxvlVZRNV5Xwhow6Mis
MMe8RKmTOZt1z1TJa3lTtiMSB8Qm8LAzHGb7KvWUn9bsUhukjOpTMMMxF7d/aZ5s/wOfWUFzOJFo
jRAsNKL92vEPUlIk4mdJMe4U3RlemydKSoDiuZlPlsVwqGX1+lCcOTCY7yu+BqpVqHW95vDjNGKQ
lxOaUB2jst6QtGwdNmfaZybY0vsfNkb/0fp6r3NLbWHsNkwYIRYojqYEOoysONO6QJhaitFIbdE/
serG78uZTRi3jxVCLKJKVF2C0JtL8ejVLrSCPtvgnbkVyOE0DPsaGgrOlJiUSDCaB4Zn3TzePH5K
5eN/6ZdeGvk+RpxLACJvYPbcL/VgegOyaX0lK5jfYg7zLSqAkzlSns/zpycHsx7+Ic1eC+R+mrRB
6WnHgX1EaBU24UXNnVfc9ovxSyfQ3ID4ctrfaf5pPrYaQhNWrIndrICYVpD2Qrk6hpDW1pf04/vP
E/goqFR0hZ4xRpqqmpZsccEHmn4TZu6rv+UEeAIRS6QSnVJ6SHMWADKSqrKeD4DmKfyhtPCvb+IN
aOYYMISL01UAdJZbEZmot0fo8njlssC/YcQ+58JxcsLIiPUnrL0e87sUMQRjWSgWq0sKYEwOMTJ9
S+Yjzfw/xaAAkqN/0O0XuReZJhqz1oNmulI0OtMOK3uvJiGQ+LGOl8W8TZrPJhjB5u0Tw1HG5ePI
+hC1sNxGie7wI2b3NCDSYYX+TC0O97m9CLVBmzmZMQN95JbeEjypdbWsa3ELDyMM9y9V0kQRSn7h
frhmNhG+aBy6u2l70poLphEVblmjEQR+rg4Nxy4xxSTVq1X4nRgDxSpD5tWmzxIz7eqSQhbLP/jL
qhnDi3ikSv0N8ZZe8jGCwtpqY7v/XZEX/I1mA+qYQL2YsUOKUS1I2RUYnkPIiCmqv7bSJv1vFszj
ZerPbQgyPCroCDpvfHOEgF2A9Sxgc8ji8mSDd9MCYmH6IkiYLL1lq92RG2I4BfIrpVsCsW8j48Ju
HL1jsvNcVwD7tX7VJH50mglHRjSjx12VeBi9mWZ4c1lVg+7SMdCeBv+0VnGjBsUYvQvE0zZ7Rpzg
5V/02UHeV6mSJqXiVrxEaifuEjC/+OiaXfjr7kJ9jIgAzgdb/HGw/cJt0hUGdMYGfWFMPIreK/9r
B7/RHTvj1V0EMxf/921lJgP+s9uup98LPJs9aW8fHXGFGlMwL+99PiU3xgQEQ9quntkMf+ieVsDi
Yc1p0AbJp0/pvMwiqH+4xbBh0ufpzGNXprTH1n3SfRwFMBll+Cw90jCzEWRoivPr/CMOi0Ba2383
R0ac48s60jB2IZ7rY9K2PaPPgI7GcExxF/YaE6zB1G3nYjPr6wvj/3GCqrU2MNUUv8jxXbwJ5qAy
SS+F0Xue4qzrJBKiZzoQYB+0MTRzN0Y4D702el6SYnxib/pKv7DwS3r40rx2KnIwdM0nGfswMbtU
RpvyXNxn3inDhiM1aXVxvlw9Jfvhs6SfkZuc50/m6gOr3IAQ4Xz3VO8bydz+oEqdu/6SYOVpUVAG
p6n/9AAyQRrilfnmSs4/bkkUxdtgP7FEJGDZUPat8AskJG3xfDdvpfwpDtO9XXANNKLATEd423Th
FTdAzuiyR6T5gXQ/tOkTgAz0wr6MFb8EHA4S2H/xgWOjHfP8hu+IOYKkHiS9IfLdUCkM5aYR79TO
P1uy02pchybvO0t9Nt3PaMMztWongFc0Ia66+m+Iilce565zUHhgectKfthPVdmO1jdFPMxwkNuF
z0KhvrzAHx0/I0p5jXR6jh9cPCvmaJHRc9fyvqemjCzXKFtY6PLpS9AqYrB9CiF08Twoqk/jExww
v/Tna7NXvFraoZc7KwAErQgvqknKqVWHRiHlI6pBk0OEFK907rem2dZkakgAic5icYZTDWe17UDw
quABQRU1tHQ8r7dzneLwbtoWRktiafTkjsJetbXP5jRZuXrEFoOc+S3uGvtd6Ox2VFl184/OxCuQ
JgHv5mdBLzcTUSh2MNfQPkrWfEtlSvtuYjtL1tHPGxytFenU1YraWvSIZXVdD034YS2MWNiiZ8jB
5qaudSYqdqYt1YT6YtxpgCLKsitL37q3eT81aj6PQ5cBdD/R9jXFz2cAkMLQyg9ff40tioqNxi8r
C+Z8tfzp2+1O542/OMuNFeIJWE/+0oFdD36ESXiXAghoUNVwqxhcl0/8DAL3xkyZg7RfIm10wqiL
xdqF6ahknPvGN50llSkiWSPt75SEVJZgfDsn97IYpcjTUSyC847kogSnOxS03lcTRQ8lGO4N2H5e
pVzupVwEvhV+yKMc90fZbUlexoocJ8a6BojqUZeQEkG+XPRGsQfi7q+Lmthn0UDfQ54akvTePgSB
HYW+/iCJP6K3t+/7u77TVqIdcE3WhWGdYybCPtoOGJ2koq6+pvLW5yEylutiQ0SRV3OprqBEqdyK
yFKyL9qNiQs3KdcgAjtBXm9gvhToZHAdOM4J/NilwU1PkDFJUElTUV/YkWt8GxqO6Vx9MiAbL0b4
cqXMviwwO9iz0XSkiFZ0sk7dJlPTz1A6DeQYE4FoO38Bk6ZUyR6P2YOsSEvqw9pzsilSLzV4XKr4
5xHFYdqMu/8HrHfpJOtd75iMqncoGbXu1X0bRsFylnUmiNec/9jh2Mlx9hSGzudSuy65Tt9Y4/+o
8V/SujfAprarqSEfgGjOgNkKeVHfb0SF1WX+Eq9C89kna1FpPUe9XzzaV/snAaY7zwFLO2TiiCSK
V/dMd7oQw3D4g0qYzpSywb6kwd1V5yN7+hiv8bLcT1jFXbyGNO82NZiI0wwC5uadSegNXmwiOUtR
gLoh4wEZ//1lee3Lw+lTvV8YPety04eeHjkf2JwY7FVkArtqUnWtTWne6x4MUcO9nqusb4VhSM1N
Vyna9/6Im93EzEcLc/g0cgkt7YRnnuU67+Sik4Eau9GWlAGkmRzwL3ceiisaz7bvfXIimp7TPC7Y
DuYK63mWVJQ0fk2mHNozUwB93FmIZdnLx4CJQJXtktZvVtOZo6N1ogjFoPmupT5XlP0yiIMr6Cmw
waZ44p8LC/l0bZbNsq9Ou/lUY5/P4+C9Xe10J27fj7kKOXdeij/gIgBAjShaAjpjtbIfCeb0O0xm
UFViLHt5UdEOj/HNyiEY6GgTbQhjpdpZnPw3riAsN4yPsZVZg2fsrV6haARqZwsOHyxdbZASEqhY
evqBft3nR7+npEEr1SAvyWIjtu5QmORunuYnQzzdMc3dtMt2KLi2ygfURTZ3gnOrHGk8jX80wJyH
g4FDnVznTPkNfE+5JTdhkdlniuAAG7L5mnxufh84R3OCxByOHidOavVwHJIOh4987Zrtvey+gXCa
3LfxkU9NiZjCsrIrs9N4l23C36QddFigUJ/sLBEOnQrd+gOrZ+dJYgywCmA89BMJGWE5k16BN01o
BN2X0npxdTgdStcqcJFnfxp0KB1NhFgd4Y8pCpGxQPbjB3l6r8/sa7eI01wt7YDp+8FGzdFnH5Kc
uwzgEV/q+95+M2JqrY71Rc7nAsEFunLqkCjbY0Cbq1QoljCU5KKh7oXKuZZHZy5m+H3vWnEhE7It
NtsvNu8yG1DMhSvLYdEnXxGnHc1Y62eK48qyYwmp12kDBrGcmEno4XrV/e+XSjJFXMHmjkX4h4Nf
WCOgli5VtUaaGu4vpbgoGMmd7LywY/25SjEdfxEzpumlwvB4Haj/6nxNgBpJR7C2w5ZLdMaF6pth
vutyJep+4v0DKNXddjYRWsIWRi2MBKESufNvRwUZZIeC5U/zRDsFw78Io+IBeat0c6bazcHvdXnm
5lPNO1ZU2RiTvcDHzyTvK8P5MWowqCDbGTfJsLuxPBpC+C3EPGjmKpxXv8bYrLPI/0OKUj+5b2uM
S8Af8bn6u8W19VuzlOU8NluKuShAyMUXnS7hwmNyayTIL8C8vbRbeI+6ROVO8t10KqL+f7w7uPCG
w0mEF9zkqAvDPZOLle6XIBgDsJNDUrUdPCSy8JTV2a2Qn0+iW3yR3rmsCpO5SfWvNswVTsHgIKRT
q3QsS2dekka6ui9jgsy8o0m1F37EjKhxmLFjqf0fcAc1nm+SSsEmMFpdboG6xRIDLVGPhDk9bYBw
L80+TYg8Fm90BSeqslpA1SYGeBxohNFvqZyXXkwdHMtzdwmiFHjbo2yMZcFHBqDkVWdiseqFO3C1
qC+tS/ThLpF1CLEQQFKSwDgbh/8QDv20zW4aX6EbhFnR6cxhqUS6x6odBXB4j7nwnO0Rg9Q+8XAF
k5dfu7a1RLxB049jyV+kzBgIecweHU2so8/GVeuoch78DdzOuY7igcP/T4gBHB56T5zJ/sdZUxuw
0LO/PANmSDGA0PUaUT2peOkGF0CCatQZ6b6jibgVfy1FN4XYf+1Ab19PTbu6C8VDYng1zhv5fCD/
Xv3IGt3jAJZsU1ie38Co7P4zOwWOAY+4DujFO/5wpPY061ya9y3ViVv2BNwgo/jHng7f1Hw17Qhc
EqR3dqV+cUxy6TteBFmufQEIsAW/OMenSlvwyRfmR1uyVfd11vQ/e1KxdEhCNq0DeUu7BlhTMumk
WJTpxS/rmOmp03/U45uM6Xy1zJjmatGfK7e/M6nhLpgMSnHYmvJSKRq6WFZDDeOHiPHchr/Km5NY
GrMlubMlA14eqLsdphZshGgd55tZwZhajxg/sDkxK/I0a91KbDZagHAGXtlrBelrL98dfWBQqyFL
An3EIf6J4alcwOoE323xjYteXm4s95VTEA69M+5+c1T9dSR1OUiLVZ/ckG9121Ua3Nzl41RUu+Uc
0Nz2Oy0xA9cCUl92zZOxaY1eIBIeZI3liubcut13ZrkP4YG7h0fvH9QJ58SN6zPZBfCEdEUgRxIX
72yIyoHx/jXhTP0Ek4iN24Qh+Dw7aiRoXh9WGaA2Dwz5AaLeBdVSE4QoYJ7NKbDObm/AKCtkCf8W
nRG/IpMaE/yF2aYhfc56f7sd5LG3SbbS8gSzMOa7EW2c0kySfM8j5dtPp+8JAzfwTBDwjWioCYiw
ZjFJEwlLSxkZ2O3V6If+QWipMcXKR6/QcFvFUX52N6yn92X/YlkxqwvTDrGrAl1rh3pcrWhAeVc8
8e813SSmDwgyq1uka1gkYlTB0oirr9KsgFgQ4hJ+g03HNqKRySZHMvJ88sAiQPmZzz9vtFLk2+Bt
+gyn0/wgbx/Vcfd87yPA5UHcmvet7p7QkgJfZJs680nF3lxdJHIU4Ijg/0LAuo0ZbYW4KCNtgQ5b
SYjYWeO/BVQdf4XPp/bDpIDfIEP1em2pR6xrd9SGeFkcNBMOIOcFnylitjzOUAKgl9/mX3a3JeQc
7OO89WcYNpPQLnlmchlmTqDN5kpI9Gcdui4ieshK7oUkgQl/kRMrGxFkko/ftZBfr3qCPjRABy0B
AoL4VdLCo/Gf0rbQ1aqQDsEZLWtljvRbX8ADlTu3ohUPAyHM1WA5uiUTTKmRJCLJxmML8LhY6l+j
/KMFf77BHF3ehqzr7T1AtMUCZ+S/hyCB/jTdaDRYxF/vCANY+XVn+5KJ2aRwayYKDxYKS0LWjyDj
/vY3lur8rlg9qhA8tQfbYkv92kHe/xjLe5Fuu/IDnt60GL6Y1WpIqkEtdalE6rZcaEWVrdGoegj6
XIyiVRzLIeZT9/vcZQiyde6yYIFsY94+LnDAGrCVkDqGhkno9ygc7MjJ7ilDwl7jbE/HSqK8hMXy
qg8xMiC6W3TeK2UndTaakdJZvCL+IluHjsiQhoIS1R0Vb8mKQV3ntbQHNW1H0zn8ro5OklDFHSrN
F/0hKtGpe6ASC4KLT5oL6h1XKAOCBAEAkxOhKxtJfFki4paLg8NNBtQqVcVSmDgB2A4C2Zdi2/w6
mmIhDPDhlOZ8QS8mqkZnIVfftY/k5hwj/voJD6n+Fz6gTXiXYZvR8lU3sNPSN8/gmnTMu8bS6eT6
91EO1joZRidvXN5NTZX+5Vc9LO6tjuiV8bst6gezI8SJgYxCe9QvmwJXsGHn/Lq3DB70AS4W6CCB
xOHkmejmo2ShPtgXvULJTBk3olIyI8M4CG762rmj2vxb84+fWytCwzP6HGf2J8RoRFo4eua10g+2
K4+tIpvhxIfZjGuUp4Zupi/LsfPRS5DWqKRVnkFiQ2gfNxHM2PvtA7Y5l5hAHoJ1ySqBOF6601Dw
evRBWkrimb6N4cxcxPotqDGZeTDn3E4Q0H9AdHKq03F3+Wq0tc8Yu785zddoa9E5kGzxiknmtg4r
BPeGAjvSUrILYx12hBlexrcXNBi3QDx2H3WTysEbstkhaFJZTEFQn8HDwZA2gskTZLXZIfgntvvz
PdpKaDaj8pXJkamPLsx0vbtFGVn00UDR1KcHTmzk4jrxL631kGOc+jwsT899M9+14js8iXGleS5t
HiLf0xayjg/iN9/KVetJdV9397BvzCQObOz2XGx7gHJcA6QRmbUIb8MKw3Lk7/+nhW7UfCdINkVC
qgsbG97iRvU6AxdR86Emhg+nFJL5gKoLYrTI46zBZUt+egNU8pMNZESUr8VOTrSCPGM26lo905Ul
+3PzKYj0y0T5BZUq6lDOW+V9nTmkL70nMfmyWNaEaJeFrYprUg1YiR8FwiM6OaHYhO2NwcFryNQr
eRbHNbrz/AL1E+bdQM0Qt0cHREoYtyi/5Vt1TFk/Yei4dJTipSAJ+cIBanBQjfU/NbFkn0sFBkVG
u6rr10V8y0HXkImpknQ50wBiikZnO/tR1L+KyrTq2XD5XUojNBCixj/H1M5IVHqQ6J3hB7ASwSz6
NOQbGl2VDhaY9/GyUqP6OKYwOgXtpLW93VJPGLSKflJoF3sDdbF+jOVt9MCLscSJ9KdOUKGD4xnE
66XMIgeJQSHHHDQmXqaBww5mPjNNRppORGWoGDftWM2lXQun8eJi98/+5L5LHRJDVlpCndzDg7QF
C9N1/XuaY+91A39LT1fCNp6NHdfEOEtpiCEKBaAqFOG4Jp1JiRhZVevX9AKThMnrveFOWgDdIEIL
XWAaSMmUhlF0ceZRSsTBIV2MJ/Ziqszht7f84UpgvxlQ/sO+QRJuI/fgrQY6NIh4/4Qv2E+SCCxL
YOeV9ygQR+r+BaVdWskmKK7pRSYNxe7s9h/ppTlgY6k7rzQ/cPIi9RxFzJBN5gGr0qMNcrNoubud
7Va7AR0nBUnllNQ1WWQxIvlQIfAqVptfCPlblcgJ4vULwdKSRq4i3CxKzoZUErbT7ENvIbbpo7dV
yxr5Ho8aju4NmRc34ISEZf3aZ5j3PsOjyfxjjSioy6UvPl9xqzsISwCUifaSh4nre0pPF9sJ9jRV
LIPd/EVaW1QvVdKq/3LFIxIt8niITGegatCJtSwhk/o0OGFaLImEbeUhFxQ7tkgJcHiG9pYYxQqX
PzxblkEl70lkJJeQKO5uIuS8w/TAyedPv3N1NUe+B3hkqZ+uNQTGDL795RHdmcr3jv8eNOH8A50M
ew6L0MErVHUAS4rj+jlPH7M9Jc2ic49Ga2D3KS85A1gBQYN2YAUyHI49ozpm3RF8ipVDG37VbWsA
RkiRxq+TOXMFTX7SPVeplVnIvXa3V3wnULnYYUTKNGT/VqmyJMTDgn4eLC0WC1yaUpPuyxIURSu+
rrSA7d1eZB59ALrXonZmj86KiQBuGkINO9KC04CYG14qe57CplLir1zfdYFPiEmWOeR7O7WzxkN9
tTuc67qELwsb4GOp+YgSWnbISvdRilqqtXxnONQ3UARyTvfh0T7dQ1Wq6xBvH1+pSYhmJj6Csmek
Gij6jqi63aHp6s0zVAgmH+KxtOOKf5b3n6SDRjLL+PqJpUNSx+jxqhItC9Zm2Yp4/2+/tYhH554Q
z5buTaHnkWHevSShzRpNbI/+ubRaxqvvhO+hRGae1Cyc3jwKM+qY8oUdakNh1kbRF1qsNwgW3bh4
Eln403B4Kag73wlAcqkJa2B0OJOw8BRWCZbBRJpw/0kZeo+H7GuO4CSlR9Y06Gsi0oTMRx/TSLFC
/nZpIWHeNmOXVxWjcl2rhDoCkUYgXOomRClD/Be5e4GU2+neLRei3bZd+nkVQcJS9Qdkh80haDRM
SczNoKIoR0+Pqw1E3YCNabxZk27lMB5z1R4XDDhfLiP1p2mLtw5ikum1gyZlK2njDWsgzoEnK2Ya
zKyUlARI2h++57KZ68JM31FSUzDHdStm/rBiQ+TKGsQoH8MjRQU5qRAqC7NIMYih8YnM27zkY4CX
YMFjCX2MqOT+U0wQwBnflvlF9/VjkDjkg26zg8S6vJBB9J6TvkwXlbASGGGuhNQoFnmLpV9WG6fq
TB+3n3pWy8kMDHd37vUfymgbcTEiSxtC/o8bhHXk6KBQ/x4w6H25YfJ6yHH+t23kneovmFeDsAJd
etef52I1MSkHkl4dQPrnyXiSGm3wfLAzIC+nZonqio3Tz4l2MHwFl6r9t8UJ0mNYRfjh9dtXw2Ln
C+7GW173+yo5Lw82RcuQC9hgpTZKyMrJZ6FBAmox48vonpsHvfqotXfPHlga7BZPzuEvoIX1ZCfa
8Vx4oAcZgsYg4BCt753Z4c6dFKl0XB8YRMZz3TnGRrpZHUQPEznPhHaAyBA1Nc7aaGBLmTRaD5sJ
+DYt0xwn8CrS5TogrtbD7DGVzVv7snwB5hsevCMO7U+5USn3yxn96ftxbJEB/f/oZbpQMpSkAuAt
qXIS+9LPE2wBJ+Vr1zsrJoqxdU1ojxFdHwv28RCqpbBpMbIBZMoEV0AyQRG0kuhNLanmLu6D0v52
7En3KsMBnGcJ9YTWTKBXgn9MWwTSN8CXSqh2e415c9sx2OG5ydS1W4pJO1qMPLnAmp+EQ0+YMqnI
a4QTil2Y9cudIlkAuU1YZL3yJxetHIa9bQSC7atMI05RwEKVhoreuEwAHDvtdtsucvNJc9C0KrwP
aRlw2+wN+FUlNMiY/sues0/DShMmrICORRKckJHoXn105wdxRh+CfA4gQO0YgKNIzWjgVKiKZ6bi
yWAwJJjs5O9sohDXWTaDwqj2YGIZwsgwjsyhUxyOB+NFzqoH2EBMEp3c2TKaKyhUsF/EfmB6A8XL
NSoz32y3cSQcBHHMOiZZjxleZP93IwGr4FchQ/SD21p9Y2ulf+Mm5txjeABTUm0IcMtOPLOaeqQD
nFEnODnutHrpEKQ6pXdTCcpvzFiHDTaN90O91BbIe3g+Dos6W7fjJD6GQOMViDwU8EnRGoj+2qcN
ejbLvvgZcAToE3IG8fGWFcM1dkMfocgSlAcPPvCEfI4Oe+/bH71zXxllMXl1kPZvoiy55jBQV5dy
30XAdrjylAhuMRIhRuOFsN0CygMiL0lQrp8NpIbA3+TSwxyWo8ThadgIzux6y3QBD5uLQfMXgr5Z
5G3xIQ4kDJTiQyLUBVUgzsY2DnSPWrfQU/3GPL3kolYDU9WbWulWA27ocUGt1WnCGz3FGRUdaoTN
cQVk0CRvsjr8yvnO+djWcZfQtQLiu/x4/h28omKzRmq/kzloa59tFCNZL4QGE8sWGVN7T5SVC6jU
2zSEqWeSlNl7gWlT7wRLeh7x8Ce6RqrHf6zDYIyKgzR0ouw7fti5BA/aTercE4hc3+6sUOVITnGF
++hrgLD02Th4NRx3CKewnvr5eX2RNelA/rKZrWNWWlw3YxJjgPBHnSkTgyXfO0hib142udEw3ZwC
sdruvHGRfQlKov0dyupm1ksLvSES+7CxOJfvwgcIrpED28efOyuB4x3Rex0Esi0IqItTza2iPW68
PE9+udpumzMyPmFA3SZlxO1z9UpTslK1zo6QHf1CgDklZLtFxlTvAUUookhuhNv90AUJGmfTXFhw
bhr+l2GKKzd11mAeuCcR55WYObViNkhPLCewbMt86U+gs3C0pTfCzvCSvVhL/p3vyU/bGBoF2T5Y
h4thCwaep+mCcFktBQBRctNciDQaKSBtGbQL+/WgFqJ5IzTSOl+2YJN/I6vRt4QecaUYEQlVpdYG
2LUuj4Egnxc+KWNqwaMA9K/KiB0CeQ14D91Zt6NQyDM01RhCT3CRwBAXs0xhe/iDn6jgi7i8EDDq
1BXnsLPs0wH1guJPGUclJLlZxUMiKgcAnFmPHHB1r+rCKGwJ/cl2kp5UfopWEjurvY6MM8ICvFhp
n2fclf90EzLoL7jF2esgie6zHzaP9yMMugRwff18ZQqqYDSCMZ7v7Bs4VLa/k3D/XgJp7V/dHOKO
YfX5U1OvBCReT9IikVYRXeLTA9K0EY2nnLxvSP0Q9gOEoQd1TMqB6wJuYtjWxRzOdVMLb0e8Z1u/
o+eaSk/CgvQrnjhtmTBS51D99kHYSrPRX3a+mMyEzs8+X2PheprD88fKBKGBnCQcJu7ad5OWqVd9
v5hSeaxcbQKidBgDHtu6G/c/Jj9F5THq9JKWYGlKMIK7ASkFyRfR3LZcV6/NbBauekyWA1fAhq4t
Nj1t05fq7MGJ8o16aAvDRdOhfzqgT/Hwsb7+8q27wYeD+qOjXur1e9DBht9ULyFOICOd+SE+M7eU
3siPWAnf/18OsvcvGp58zJ/erGswLybNZmChe4CsNDH+XJRopPoKCxU25rAY4L0Jwr0iS3sdF/Ov
8F93TbjzLEddhWiJ7fpMQpL3fpZ/dqmRv//qgHnuoBTpWMshC20nePer1DE7vXiSI7WDm/5NjQSZ
++KhjmG96s9qGHRyiDvUnuZK83Xk+laKMepY/9aPnYBUecQ5liqENY7OCh4uAigt0TxfloSMBwRS
1yX52dtUdV9I5pWBe3esvbP5LhNp70SSp7JdpjON4EshihlrMAHybz/wSiSYPqgXm1v5ZpyPtgUF
cQVBaDHSjB+bISuf11wIBOfdsrsC7/r3B/yxeeUEbC3hJDNU9x6ClWnwp9INh26O7DXyQTf7COll
YL8S0GnVw5TLhPo/ih/6B+1CEfThIY9u4ZyoXD49RQZ4KlN+hQCfnz40PU0KmwQL4KdoKz/H8JDM
IsKNiGBaDB9TI4hqiWhlpVz4oWC5bGfcpFcxNjCFI3l9xxqSkCAi+s6BAq965vbsjMiNtjvNfB5w
4GEsjx9BiXj6vr8HRns3aDT2nb6XOMFQreH3NdFgRLvGDiAyc6LkbtMBPleP46NLGVNEdwfv1I0A
qtYLTP8pX5rsEB+ocnnQFSIOR6lP0jFJJpHvf8FcFBwwCH2rQs6bjIG+eYzV3xQ3sncopUFINbvu
spyJjM45SXYIBO4G8S5/tArushTjDhGUzayw39OLJcdGM6JMSGQ3qA9VGsdx6DLmiumKXXYNZzYT
agr3oY7AwSJO274xFppIZUOtz+PLI6K5YYke2pkAAi/HXXPxNebyjeRkZBKaw6DoH9XfWC/tDl0E
Hcnr+T9pf45P8UeLrwdjAqbyj1NPUZKI4DFbZmVxx91oV30j50JcJ9++3+Jej9ajLDSXU7y/xgVC
hPvtiG16Pf1Z0hQI8KciL1Y9acL4qPnPGjovpUK9oLKg9XczPVKo88akt0iFDAGCvH4fH6NbqZuS
jZQC7vPyN6nT3GZRd1q+CN1uodg/hmKZ/KHem17GH1AFWt6qvMgS/JhKLiqU8+VXI0voiycT3548
+YGxyoQnOwANyl+tuOSEUG271j+ndvKDi9hqBAv/u9pymu+RpVyezb5DV2NUAZBbAA9CvF+CWgWl
hKjAANDjfQnc7f1Ad3aUNfz3aXWGpOW1kQdn0mpqZjH74tvvnES3pzh+mYu+sfUXiN5uvZLc3cJf
qv4fSNTJJ0xM1oiO+Y0k/bt/pja4naIityUtaQSxGsaGD6Yza5/2nlOmEAojZi5w5EXafdGuamod
E2WPA+TI3hvCKImSRsB0gh3Nz5RI1dFfPP2nm18E+QTe0dw9FM7OpfA8JzZsKPhhF0FrcVgSsJHs
OSU1kpc1RycNSIPjbJ0qx1tc1Rjrfv6BdTm+cnp1QMFlZb5C444XvWHgV5qoWiaq8xONV9+0BR5b
9o8amMV7cyfGKiuvCvxo66jQR/Z6ffJ4/dgsgaDEUuwjFA+dqPhrydOb/7Elmd8AkrLnqf2n5Kzc
EF+rzVh2E1s9E6ky3zXOApv0ZLBnXIvQYyssi++0XX5y3dfPWJnIpkD6ejIA4Y9Hd3N3HPwrd/Wk
ZL70GK2uz/M9rSua3PN3LpUG3jAjzIPwhvH2I3c7sTxSHaU3RI57Pg7H1SqbRehnkg5vWQn1mlcw
oT//muW5NjdWumJBd3hZ5AvGBc8cyQ7vqbIx4CNZqz0H5cL5egC6g5RLQ27ol1kSwJ1eP90YbyyP
wiwJeZ8WG8PnPZE+3uLEaqUtUyejjJ+tUu+en8UNeQC+vK+2sYHXKAfvAdtMY1Lpe5Dm7giy91Rl
QDEOC/EP+qyGzE/oClr3y8rpBEU0x3vTK4rDBY07DnotG3ekVr+PbIfsZvaFxXRiEX5bGh0gaaJ3
Wj3tRU/yOO8m1CSwPa6sqnO0o7kz4a4HttdtXiqlGyzxZAgEg4kvVZ+oKEZztGQu5Mra7yLrTckZ
cx3Raa0/8N9QdJ/BDt6MlXA7C2ooy1pS7yvWKvw8fQzGccS+tQMjveJw/Yt7SzY38Uig0mrd/crE
xx1MdEoRjSPS4bDRXs1Fl6esNQGP3YECV+J0GId1r1uykmzCX0v7HqXTH95gLvXKgF2WdyLyjxrg
q0wzcJNgaC+2/WfwM75EnWmgoOe7nbwCsICEkpW7TC8Zq7Mbb+lOBuWs37QtXh3dOjODdMSYH+/p
kRvUIqSnZoenu0PHPffCXTXchuziZmYelLfGdRaew2moTrdnnAT0jJyWVPirBFnB+5o9rC2a2+cI
bxyxte3fHxTJUX55zxzkN2JX5Ta0XeRJNA3w4iR3sGi8eKtFY5o48oBb5HutnIH07ski6AhfFm3L
HdttBObL/NNLPAkSZFKp3O7usaGtilHMcdhckiT8ok6n13N+XBHyV5w/OaT/RiPkfC2UkEGrvysI
Nfpw/LyqZFc2h0TOX26wZacp0BOQIQmMU1j/HUAauDgl4zyCQBV3O7HuRTg247DFGMt2XxdbJFBB
fACZyxrEB12K9yJfgDi08pJARN6fSckO4c5QuLo96ceY+HSczvreh4zlc2HdyDg780imrfDEoq7I
RcXplJGBwGp12LmhFZAGEMTkohiIqYl7929m3Yt44lb0O/YrkutbtP7EWQkJ7mRs2/mZ0Xr70tBP
il5ONVFhEMKaSuoYO8eptu7OJmoIbitiIh9h1RbsX6bMNC7eb6j4hoIrpepNYNpLAt5Y0AcDZTcu
YePa/2aGaTJYY39EIgdLf0cgkqQ2Plwkib015QVD4o+tqYROvLLDZuhL1Kt88NGyn9V0otg1BHLs
3mmTyZRo3V/XvyIdTNB/EWuv+pGAexFdVX+bFCvgteGOphSEkEqxYQlbuHdHhCV4DeOCBCMkkw0L
fnKYIhfoUTudaKQtvxCrVrL8un0m8fZXuSHN1/GGhwIv2zdWMf+vvmq6VMaPLjTkKeQqro+ZxY0G
//m15YlkxCvLtLYWu70A4Aglz/stw/EzQfX+5VkNv1sXZiBAKLeTUkcTDFmd6RmVrgixCD0iYA8t
cZH9pfkuruCFJ+zkq16/LCfP5AGi9AmG+IYbFehfA7YbWXfDEe3ZWdHQkicZSANMpHU/OZn60fRN
VBCVsn0VkzuzFWfstoTwOcBbUJ5G9m0fjm4z+kEqOB+O/KWcU4mGWqQPD78iHkRTvYxITJsvL3sq
hWKVbXC++DaRzlTxeultpBpAVxRxq0rCy8N7hVJxAGsEZlPt5pyl7pAwwbEFLYyuv1Axgi83+ov1
vFkm1y4XnN/TH11qtvrlHrcT5ILWba7uVTJ4Vc4uEkljbJzUpKvcE2wTvL7LE8qQW2yn0dyv1ATq
zrnMC+3bqQ3LFofoIAbP6LgStZnP6VLdPLovQFcemaV9OcAukD/MmSRlA5xfBFNFpvnt6EtJNkcY
3lrNjwZd1RE4qyHkQ1WkOwxAGf8zM7O8mt5ziHwaCF1LqmRCzSVs/p9NoNcL7Ezewc9dWL8EqgMu
3zLfVeazv3HB5IiuxO2RZSnO1+R5wLJGMqZxuxEQTRkvSHfLT1KSTdIHqKIKr6RnNRGM74kA7lq/
jkhDJdmWKLCYk41v+dok5cMIBT3xmzfkZlSUb8okj4rf4xpAFRa+MsanItmfgU/cNiK0TTEHfnwL
knxjVWNwmuEpzXTog+o8We0I6mN9di1b2JftGz3yav9BSj+bPbHoEGSSfW8aSKO+YIZquUnRhquS
OS7U+spBsiTNU9TrQ1wk/h0x7t25/7rv5accTr4MwMwqbBL3jRzqQ6ilvMv0NHWf8053Qf4ynfze
fqsQWa1ZQsgf+z3O8LugOxQWachKJnvVZeAnWKfTPIGlwxo7JwKy5Vwxn/ZX5rTiB0PaCsnDurxg
ZzzomN34f0niQokDeqfNog6wnJTqMuWAMYaWDt7BzMknzb6ayClg2ZejRHxAoX1n7wPX6fhUj5vi
YzL3kJtSyJ8YIpLRltJXooAsXzzkqNAUvWlmcN3GXvIUbh9PEkzcRRiHGw+C1WkPN7QuWM8eaHhV
ZPB2fvL0kGtrcxqPnEsDhwSgDxcCXY6XPcobJZAv4r2sd3VZQ/2GkCalhBhSAdjOs05N9d+ol9RG
jOiAAGyrUdORODi18dVSneFOcXP8SGjxLst/4NAYU4Gsp6uWnonRKPLZSSE/txoS3H6y4KMAU2cd
LlcIXPoW8dY1XcC17uzIP8qnV1I9gwuZmOd7FKbpeYlELcFd2hJrWmqyuRf86J69ZGOuOvfSEWWD
qtxw8kmNfsPGkj7VFMPTaHjNpiEAjCnHjLSIsJfeQEx8CSZF97RM5E0ounY165ogFaZJbaCnck0v
yQ31XBW2uGZNOQsGDpENylz7lTpKtoNtto9YBm46sN78O9vQ9760FcxKbJIxUB+ca26Rji4si2Gg
rRzsWn4t54iCYK68G6EUBM/lf1cssMuGu/Tqa/DP005iyoPmGFhmg8QL9HgsvTBPK3KbM67JvHWF
pWNLvkytmug2fyN0D7XZ9LJHJvyUM9t3XGGA5X2bfM8b3WoJGApZa1kLunbTORXX0mFrZ8h9Yj6G
qdstJd/L6SsnPNq54Q85qlSKAEUYLoBsH4Cu2mQEbsNiHWWu3nhGiOpxzq7Esfc+jMHgAJs4C3N+
FdTVF0T3fjP8sEq8GSJlZooi3H8ueNZGI/dItbHCzYvcNBCScy47tHfL7qQT5xNTtSpT8Opkrz5a
as88IqEUuI6sKY8AQNyXcSv/XYGBzSuAdz+snzAiIANypxtqKMw2479IdeVbsiwodRZn38pcPjfp
8hOGUMlGB7j8LvCMqL/1PVR0hXoEmTjw2DyzIKgHsU9jNpL7MFw1YA2YbXDP3zr8YQ7YNCrSzXnd
hfHlRyWRtT8WEgehEAR7BO2/Kq2gSGKHQIY0bz+m3y7Lg9hQ5txW8q80PUf/5wSEqBSRnXlkVPs4
uZ7l6mxouOqoltfrqTs6GnKM14/ul93HTODsc37S6XQHq0FuU6DdMfCfo/ilJWD4RnxAEVlHF7wB
Dh0uebieurRN5mrSkhFGcDJX4n/MM/ymFN9nD0qqQB9HqckgcXYDFeuGXFMcoI7UO7Jr6xo1Cq/E
KFvFhw/0P5gC6i6J9WV0BYhER56iBTKGt8CAHvJslYZ3oe02UNyvvVY7T2ev4wdbmnN5yiegZCqX
k26+jHitWjN99G2+89V5HaWfSLdk59+pQXLRRpvkKVXT5+4WmmM6PAyUAVCbrgbCXuFphJ85vrm+
VzaFUzBh8lyL9HytW/Spb6ZkP6dVrk2QS/7t/SmqJ1iRaWDuUYzf6pMysn/1N92FCQkEQJKaov+8
FXs2b4nEjcB1JaXioswSkh9OF2neeBvdxgzCcq1uwZHVg3dViyFW8dCvj/xEh3icOHxDRY9515e8
ttaMg+ZaBB+UpYc9rjxhjuF5TmEs1gD9QgSSBn0hJliy5IAAZopLFiezwoVcq5+T1HOzwsUNsQ55
mjNATIOENrmC3Osu89hl4AXCJpxBsh2FzuR6TqVh1ukRubjb40qFQdDio2gF8u6elGZuXwraknKH
wAr3cd3wkJfCUN6UxHVLMRRIFwPTcAFB5OdyMYxPYi0seApCJY+xrguS4SBputJacw+Le+/qXMqt
fZxNTRb8AdN4sZKPPUYVOYcAETFpGtHdypi01rTvXXGq+YvAq4vLER5X9+OUn7UmwfkTveuZ3Jll
Pmcvho1smda/5Vuhcznzz5IjNQMnGYJtkvbjOZ27BgdErH3f4zwEbzCQTIyGiTd8Ik4XMLjsvnlh
22oerVxzYyemS0NK/K791QXut23u7q+BR2p0oR+uY9LbxOPpa/f/XZFDvXCJa/lDQ9TRwnSqWEWV
xg/ypYtmyFFAgeBm1w7WN/xpVXRjgvoQG9bCKts1PCdYKSgplwcg9EA7rALEH3lmKEm2QKY8MfAW
XVIrAU37Bc0hDYjXE1YWkZAhI6vRXud63P47X0BiTaKXAgXZHW2EIzwF+h6ox0eI815+5G2kNwp/
FlpqDTSMS2VPtz8pIY4j7skz71SYm8eLAkmFaMLKyJQAQqQVJKEKzP8iJey863e2HmmgccIu8Jaf
2SxW5/kQCzLL4t6Frlro/+Xoleho09kWM3lvpvPmX8QPREw0M8BvjgmQGIhWIv70nNaKPrgQMEfw
dednVGYo1GkfkIXp7tCmhdglMaRRGbCcMhwg03R23CYjdW/1eml5E+vh7EKDpXiX0vzeSYe5OxwV
ZzKyKDfRG1sqeUAzajGdbcPbjeFE85AlcYBduMNX728TOcX2QAuvNClbq5vYiXm76mzPmyNtZrjO
tNTm81g4NaydlTus8hQl5zyOXNA1dL3Qva1XYDHUf/6e/CxByCggBxmLnkfb6ZfkZ+VAR9hel+Gt
A1uwP6KEDxVbcQUpty368EEXAkco6FxpbihHouDbAEHfW9SY9jwXbWu+DtgQ7w5KeNiLFqaLUT62
saoCRPNV7DtGqMp1u5vhJCCDAHOQBdirYTSf/zKN1XsxjX5YygPiecdxiYsCWcadxEzP87JBDFRi
1p7EtrH2ss3j15QVH51WMCmVkkPEHQ44kmIWR43z6LagtJgcInEKMa6/FeEJPTaBurRhIOU76hJP
RDdA0oBBSlz8mrbt0kE6YbhWzPTpxmwvJ7n49Wu6pMono8Dmd1T5X4+L453/FHSNP2NdyAyL3GLg
6XLiPMcYyDG10Wq1fqVcFZ8eFIGpJDmJs3b0Lb+Ad8AUtL3MOXSfNMqar3G28QdfwK9T7mdjUaw9
850ioE+pTbg2ZJZSSA6HQNlbdBGOMBn2NLhL/f9ulKlTGvtI0llnGDUuX70+9iVob41eCY2semRN
QxdODlgm38g4Sfo/2MypjVCki0r2ok4yxt/NC6XMBi4GD4gVCtbDIMfTNgvDDhBHrxlfCUY27KHe
hb/4MF+HYX2ly+aW5VFejTPbpYIg4q4ZY0+02XM1Zt52NnmpMD+WsIIfR0GUNdmRy51rkaDJ4rvj
X7KCUTp+nwsNeUTVwjM7lC49K1KNoLd92DFWT1p7AQBeDYU999AgJo2O25dRdSrbsaUAvii7juGS
308audYuNLL7pS7mLJNDwY96L0GxjBqFEhz8IXEBhzjVV/3NCjMnf5pHPeqEjBcGrBHmGOiki0ao
OdcvQJQ6yeVkBOgtY0uZgcqYkj0NozVvxB7PotOkMHgIo1eqyj5A79J45atosK74uS5FRWit5pIi
Nwf+urqWQ7s8/3B4N9QQxOjdU4dmM7ZmZz+BTxCF7VuN2B4936jTBJVR+O3Xt+qOmYTVFAfGcUMP
pFaOPf18WhrQv5ZUDizVv/Nyzj+hUp6Myu1fJ7sVD4PCERQwFrHjEcwJk62n7WlCXiJCE4L6+9RC
qzlfu/fhN+fE+G6ePtplLf7PCwLkdYnAum1RLPUo57w3G7BOtkqMwRQX1baxGaWhESw6sZOlnmR9
T2KDb6PPLeHJQ63wwxD9DBRuwb0T2SS6v5JnqKXl3TrQOsSdww7/r7RTUnqoUE9E5eYv1M+ruEK3
oOinqOwSe55sZN/kN9YL4aVQQ0QkHfEVIqb6QckYZ4IB3oqExjlSuM7SmeW5mGqTSP3V7iWexqbw
xogKoTU48n2LzNdvqfwY6b3ldznHYKpzI3LMhNqTZeh9mvRreIk6yxd+YWSIEHl89JZbkk5OeEEP
WtsUrprK79Zx31f4OATgcjl6ERZrsBZO8XAUZ1oMqZ/2W1cJkjA0uHVsRamCpjD6ulYk5SzgSb0V
/RFHgCLXX4sbNJnSbmicT7vJjsSoNHpfHu/f6eJeKaWfaJ9LcIAd9aBNfzm+5E15R4N2iW+zvzD/
zwsvQ8GRzs36kDnNsHRj2gKO7mod73NUpb+3+e87R/Ak0KocotIHtULKFTF1k3JkHeyawCeJNa2p
qhJqyMwa/JpuOV5zE3UKaOcXieYwjs88sv+8jXnw8lZTp44MQ97z98ZJu1mWmuXHPVgMKUE7YNQG
sb6qPE6RkJ2byS13IQ7mEMsLhZTbrk4UE3iCW/cw1wqrAkW1p2PEjN2zYVgW6jzB2KZeRGPCIJeB
m9OOMXdgdsqGpkLTEqtPqVR6HltBCHStllzZypJ+MZx6J428dTF3ASibvUr2N7wKa0rXq9De9j2k
Q2Z0P3ymdks71/Bm/bwgPOwbFhzavSNXAuuu+yA8+snFzxj4YA+G2367eXm9PkiyUGYWIDcIjdFH
HxqNgjMiUuK/ZSAGRlaYDTLieYUoah1bvs6Ub9TmV6ic6/Mw/6jQdGXMH6OGGzVqdKyMXRkjsPs1
+gxOFU9WTUCUDOy0ERmeMwD5XATjOpW2PmyeBUot6OwvGm6gDyHHnUIV0FLemrYPrCygS1RVwU0a
wwiJd6OHwM6YQ/Hu+huNPX8o0anna+WjgDQbp98KeZAOApx4vl/gRYN7lweQ0Kt4ujQCvAI7P0Mo
IiqzMsneHru1YQkJLyV1KIMaB/Bc3IvlmcoQFd+n4+nLRFG/0rMn4Cfx6K1YShZP2XkV4ELm3HcQ
PuZwmOpVrYeKgokq/GzqMA3/gXnOraZ7MgFlSU1064J6bGiCRyPtG/6wcZHj8tCCrFPr7ie+UNae
nFxewRET5MeRUupipzcHthQ38vb1rc9r/ijJE9EEykh5M/S6BiigI3S0eisJ4pUu/he7KyKgOF5T
TRmEus8lja51YoHsrzCxRm3MFjXSsJPjj6LNzFBUE7cZdn616YHCSkI9cW+9FjKWR6D2CxKZ0JP1
Y4v0IrrMGRIgG6ARyPqmJs/lBXB8vvUwGarS8BO0lWjQcwLQ1ZLDJ3Vh4eEOpV0LFQmaeojRuBYR
GQc3BE9JDqsUMRkTAv3yOE37T3qQ2qa2nXCU0JrRsIxTRrwz3WftKiDWpkalbpIFLnUCXwFPq9xq
IxdasQluDtb4odNl/j1N0tnckD4/Bsi1GWq0UUgT2V/IrPW9+5fTc4WKMFt3BGBvlTeza/xBKT6S
Mm31P4YUOOS9xeJh4UX17s3Wt6dICTYcdm+vzNsICZdKjzZIQ1tuwfCpfBALTDF60YrXeO7UI3i7
RgpEolIFC7J19rZaSviefYv4PYPrDvq5BsEYK3RC5dX9YibjV1eYl6yepZVUzaOOEJ0K2UnPw+KG
5nVW5VsdByNueMX7rfKVU3F5yIJ0DFISlhgjBk5IHCfwc3jpCee/S+NjLoSXVlPtmYa5jXS65fAb
qklS+9daoVgLbxC237QHr/2QlPlHuBCFnGmPxtn1HULPt3ScoYLgMATylFClhjZCuYSM/yGMTqJY
CZbg00SCFnlmhDRB8tUjl4BfFl3OqCkITxmqgUwtg/Mbv1vEZCq2w31/B4kFs5fEsFsUMkcGtQSH
XMPRTDUabikfD9Q8rwT1v4a+k6/S+lj2EffdvY+cpOo1BideGmD0u5jTeVJHv9lIbUb6nW2w0GkI
Mudb9R4jCZBu3oDCG6EtyFvIVBk3K+TcZ+2wx40VFfO9qXrIhyBcgwtTGy4SdfIDF3uQu7F/pJVu
DiIGmZZ389A+/3kBPH46VQGFETaN9EigWBpNo8xfPUrhQXO7QLokKEWPSmgHonsnCRDp3Omj71w6
+TehPf6w9RYFdmoCZtsNSK9TgX9lup509TJK+k3uonet9WSzgL1jrszXAhWkgciuV7v563tYXi2z
fYe+vf6VhF+LKv0eju8XhkZSfAZKq6SCG44vn39zJKsN29ueo0PGb/9iLf1QTbRrc8Z0DCnasLKD
WgC9Y7Mf3qimzxgzPFSTOw53/fDeUxmDyCMt0dvHvFMqlma5OarmU5UTwm9f7bkjMrtbXka0jLAr
09LMtkbH38HhSjs2T5PW530xF6qQzuOgjIF+sDRzqreKWXNBkJroM5tyIMbHEFD7dzPsIEWM9Z/F
CtHIBUJpwrI8sF4/gm/qTDnG8nyZHb0p8/uPwW0pndEwmQIWD3ep5Cyk6Zmo8Apak7QLZA4j/GZd
+fFMmfu/KSIWYgcO2UQBtQ5cj14d6dC/YxeS5x1AbGWRPGLPyLea0LA3yr2KfR14fhB2xgbxWlmf
PPE5UhOVI3vV0iC2ab/dZPt0wCJLZ+kYBQl2Bkz16+TqOkCAQ8WXB5xyndlzvsJ5b1OV4rmLQ+FT
Acv75qt1qwSpeiVtERoKD2qmx7I0+q62yI5JzsIQvVPGF+D6wmqKkfsD8u7aooGiTbIesNbE0INU
2Y9ZRH/cs9YEipLpEKCOgcsn4l2LS1Z1nnUf0PNVO3/JugWkAApRJxbAO2DntRk40MpUakzf1OUZ
EyETAG6+s16GxmmnmdKIHxRSnWEOZJ694s1/7cQGLDNIo0aqOY7GUbBSAofuEKCAeQxkLYGlZn2G
3oe2s7ZOraZNaJ2Rm7DxfqwZ74p2RSpFNAumTh0ndLqyotkIcmXVvfCgM2rG55bc3v5ninl+lZ7z
YYoaOaAqeiParXe7cMPDu5tgGYIAOCUk64TKWXegBcj/aKHyKrbbMsY6JLu43JeoFYv3zFQZmZRE
e1rbyqwIkxGqN3QYatJSc6dIiLajv78lJu1Gr7HDPTHrFRcCz51UrGLOWQbL/w2NfkJzUD3n90QP
wa8J+PCpYkDrcVS5jyHc6v4hoCev920HwfnATfH7uuLS7lTnzQsjNIPOapk6bBdn7OMGZochtHY8
CFUTPLfsY5CPs9XSTVTjRX3suSpINVLyNtVClBzUN4VxPYYQcMSBvO7HabBzcvUcbdmr08j/ogrh
mAoNBVho4UXFIrq5OUqGqdECqFZzGnSmld6SkwRBpn0Zcd1oFkMDilBVzBiGk1yqBkQXRraalfTm
1K6FtvBlsW/balJzihiWh/A564pvhgdM8iKy1ElDBaAjzus/VMdRK0Fs7DRCZlYOvZ1NwGxngTE9
kf7zdbrTO2S014Ka13J9L+EW16Aai9+o8ZzIneDHPCPx6BehQMADrOLfa0rM8MQHNzmlAd7Ik/l6
ZFYoUKFW5riVtY4yHAB+1d9CtpYfSJfzrAi/7WhFljwDRSBpAsiYkQjce1RDKKED/jQVLB3N12x7
Nq6gAo1/XpmdR+HLsRJmUG12pEGljSFAtDH1bwhShHGNw0uMx0xW5FZiMzGWYC1zxwtpQWAHcanU
j72SfvwrUE6dAf3iZtk/Cf+D5WC7bJgPab2TxNe0E8qKNVDXxlLGJcKJLMuxg8fVxBjO4mMm3h77
mVnpQawtM8+MwtJqt9dYTJNAxeLbGZ1H5FlMljbAEEp7TzQ9APxyKPW34/YKkANp7BubaVWJLejh
rWNGjFB9p7xIJ1/9nM7x0fHojVtJBEdwKQ4rgbnNtWHFo5uOaFhXOjIArBgTLU5/P6z/kHtRRo8t
9DjIE2VVqbJTchXf/f1SsZrmwM39lZGHftPq3I/c2lXtISCzqYe6ySpxwYg0sCv+JqueHrXJsdNj
bWD8a0hUO2o2/lL4DbDa73eIKlkdvGRWrvE+M5ieQUZagmN5C4ghtHgfGPFFTKJJ4rYImMI5fjgd
ke3m2F//9YMJgeXxA+6kjh/dbW9uqwU4M40LA6gchGCSj6Yp/4vCQaaaMyEfZeX0R+9zckMWB1v4
T8+RmWQfo/D4o7Nv5bXbi2d7+qKav2Bq1pBmY7VRXFe6mf5wIr1awPQmts9zjUozpGSmJ8zzJNpt
pmr6oZm9r1mCeMUJOlPIAqOCOkt1Sc689VnWCsj5OHwai5QXAekW5T578N6LcBp+gYE7VrKHLA24
OJlLcbgvt4kPWfM60zE4GHGTPWDTmmRMxSg0ZXdLzOOX2zZwAxA2H7w8GMqqO8ouwYNI2Ak9k0Wo
jOQfNIjukwlFDtsVdNTb0X9iyQZJc8lVke9xMXNSFeNmMPS1mTXIWUYFwEBWOWFax4WQ9CMcy/eW
3ZzK0LhxAytt8/Eq3avyA14dzgeQ/GhMMN+YSndRvjSql+5CvGrMLMUOctefXxqd7Z7YZSgexACm
ZxZ2iooHyTEorGdXJrpQfQ7BQjUCllFxaFsOBud2mFcNvWMhcZzDmBs/G8B0UujkSlbGDM6FgRcq
CCN7Ff0/VIzt4455GHec6W9OKgGmm6E1BEUjSw3RNyVS8VHgNq8PWUTFKsyqfrXsjlBpUDp0bPdI
1wmJ3hajqvnaJFDdFfXVz7yjrbpyFqBb/QxN/GTuU1G//dgF1U94tishZSyvOl9rHLlF1oe2KOTy
oZnweQCCkvTXTcno2sEH2uTxWCVIViw4rXjXb9BnEYee0aJwbUveCgHM3EqVxP3+Yjli5Vh7JOwK
veSA7UHSBYoDvGBTZmmGhef2+PG0sc3nIvElf36mWeP0+ux2KNTNIBiF/Ekkf+JPg83RHz15nxzT
V8DZVGRpPG+vbFw3BKPxEaBdFDyEM9J5qvjfxb8ZpmuapalNUGYK4OAo/H63Pa+ecOCO3A2o2r6U
qdI0kD27HSpcKCJ3WH/Ax92pFaonH9wd+uCFJutcthgM5oi3BKTSG5pWTLM+0iyHc61tqPE4Qg0S
hXNPsNB3oHs+Ra0B1N8leUvOKScE+dBy5esJKtyHA3bU/1C5XQuNrq/lLDMEsSvYZ3gdiIygYibD
EXirRIDEJz+h+/8q68AONjCg+0zTikxrCEEOuzlP2/rGlaBpkGwIei4+x8CZYVue8exYga1l2iP8
Q2KQstFa2j4EnXisuw/CRDD9y3EfvxoHqsDqzQnrrilx4+pKyTnxNpfIQjLsluQfd1KM2j6DxTWF
k5TR/FR1KPt/ALXuaOIaJuAp6BZoUw9zr7SUVsxnDrffWvE6pLLbkCWonPRxAwAXLDd5Lgiw0Wyf
wuzjNG5+cwqXuuqSt9isdMhGW0qiQT1ZcHu++pJs95NjtB7GCsZ68gzYV0S1Y5G/8kxw/5Fl3iou
3/k6YYBY3/GU/kjyU15QyewCPjk+iPSJcyci/TWuQFRQeiAczuQuyVv74gO6kUcVKvxmu6Uy5+d3
fUaEdeX/EBrW3QXYeUaeEJouzxwPr3lsJcBNw+hm9AqX37Ym5C1NF6JPlpDN/+RDohZV3pwJlbuw
XxsmQ71sIUddwZRDpqxW1Y/p8GE/UsdCdAu7ZKmBVixWezBXpdl3eVy0KNZ+cW8HV/H/nqxrNldJ
/tlYQNWRrjl6U1+tNmLhX3IEzXFP6lxirgh6ZIDRHCxl/cz99qq0/YqftMUbzaKdJDtLTR4j8FHg
tXIv/AOStEQ3Mcp0XTmwn4alVgcUS8ioqKDBJV5x3LEYJmXHjkZChJuz3lQsQ0ZIN0lTG4r1zKYD
X6bLg8umDcoATWYNGPPcmsp7rqexenaClc6d9B93viL7NcHgS65UbQcPiUMIMtBqqWPxcnImN4ff
2puuD462fpj/x3n8VOTwoBkWvXQMGy045XHmJiiXFGi+HEDQufWHSYEMFlE6GT/xm6qgfoytKawu
tjCQbkCcRJ4y4+fiOn9kxjo9Qe9xOxNktQK6ZPH8YbuD3vrnYN6L1RfCFEka4QXI6vWwSQEpd0h/
oN/GVLMJs1JRN/xdtjJSHjQLUWWhd8RXAOv29tSuhKM/0FPT5TQcbZQbqRTcWFjnxnYNqS02HWsv
R9OJnRNRJSjQ+DYWx7M4ytFRGHB+wRVe+5zJicYAX8+dJlEM0HGKEA8TDUToICb5T+8KcNWHYlXN
uodyNqvEBEmNGjEVeLafEv40Pgea47xp9t4S7cMDdLGa+Lw8eAbPgA+anS1synYpR6bAvwxRwcaR
1fu5I6hrsVcZ69YKwD3YQXugAMxHOE/O1uxlO28+t/zPF9pbsBWmdhaq3Fkj1nClO2QUyqPRD2GB
Z+WgX+oNy8rp2AUEvcJc40OnQkUeO340s+QL8Y6sCCT0HTzie+X+diqoN6X6PqWeTqOi4lMDoDRe
7mdPHTcSOn6vjQSlxdd+wlcdE14vSKUtVZ3AaMImdN1SNHonoXOLaobx6ofcsUe4dP3HuG//MhD9
sw0HFOtIUmHHIFsO6Ud02TxDAiQLUjXv0dC//qIB8LAum+HKOvm1otvDS1unPB78q2swO9O/8Eu+
z2H8tkIuZou/YykOd4NS0yJjDwutpSG1W0d/gXStYZz+uxqSVUYSeBPY9StiOVsFneCauKfv9pG/
brpUNOP4hWTa03XVrfDp3XEmD+jKQOlYCjrGsrjiz5UjH39a88uEN/3lsLeEvqUA6B+dB7ubKSfD
FGIMV/Awk2WeSMdpEPayX1DHScpetq4gaojt8CalIc7/xNr2Av8VFp4CHb4Qmj+H81lohHUwmj8+
qC6L9aiD2aPf6ySfu9tXm8H7NWH+8jKiOAWHFDRkaXsRZXVi2V+Mtm7qjBK7q44kRFXC8qfpwg1B
LXiJWptlTAE090mVfzkG1PnYDOYLLY465tl8wLDvWKL0Fzyo9noIQkPCDhiVDGtPijeFICOOIi6b
wxCLMc/ZVXMa98MW/LTHrd4ROTc5BWyd5wzVti5F0HShxmMBSbcWNVRyLq1/gmXgPjY75H0rrL5S
WQq1LtFBYXVQxw7Uv3uBC+Pe9vRflBhThier1CJZN28l/CfkGcb58OFD8QtFWnQuqFvbxMeqd9Hv
RQIARX3KgUJFR1kIFqwnH/86Sc4Pu9g/PdlmFarTZQ0WB7/IsCH6E0K0Wp1MDgSYzTdWP3mI3X1K
mxChEvcnn1KtqlpaswqMv99ni2idfduq+QIpZp1ypwVuAJQEXDBmkeDaBbNF8t25ZvD00xs9QCOl
9bK512Cu0R3lpTkKuFAfI/9zqmzKLga0+2xA15sMt728855ng173mawj5kz1+omWmm4wZsCSFN3v
l561ucW5a9W4Ff+iEJPk9DbAkhcIUBtlPzZX2bOWny2Tg5Ai0rWwEWhO6huZtQxSz7iygyVVR6Cq
Gkq+TR/4V2UlwJaPvWRsRz5Be5V8PfIH3yMG8uiJq0fKZ0lvm39rXBDXZJVbM2v/Hdwd8JmUh/o9
YqQLTK2ho9dnMXd7KILADVI6z6UgVPPJjvBkJw7lP47mHs7x9t6lIYvZOgGJW+pxRkH10jL7XG7H
bvJJiaNoEz6zvt2A48lgUh/NFwi/tb+59gkbhIv+uOv/ku2Z5+4w3MnvnAzUnxyrsIM4lJkqYMyX
X5O2QK9i7VsHNrRPwVXUucCgODYnCZJdwsT6TotOPHwQ9o8+ggYv/ufmGCSBu7YMCAd9waDqrBZm
CWpXi4hW8fuZOKiHOzYDuzTKG3iNJ5KfB0KDqYw5CAABJZaFfmrYNhdX46IJKYeJ0Buielb0diLu
/CdtV+SKYJMHm5Yfn6TD7wTWGkKc/qClOehKPKRmnGwtp3C4yKKlXqzU92/a93xioECgmGLl/Nkg
s5xYoOJMlUsYxqHdkkqha4SRShh5Fn+JNKi1ZRL4Co9zCadIVG4DnGBiea+NkgqgYNtvy2H0rt+0
P7MteXCWJ9ZXZcEZJh1Zn7IWDbPnZgfMxorrRjkGEAUT7S42Yo9iJvy1Yk3C5pLGOEDjX0pjBvoK
1NnU9WDEN2qHrLdOn7Q5EaJKb4M0+LxATDLFY/Rm/XkzigmIc5K3qfDqrPFai2a68tiDPtTalErs
CeI+IJ6bMLpu5uUC1mfAJF0uzcqgl0p4HtG9TNq/MkniFMFP+6Su2azkNQ35oEk/8N4oer3x3KDU
kk14NGObuJAb18/QIiHqU4CRaUVH6UfaCkGrVtIc0w58eeF1ScdFU5V2PhL5zKOQW/lIa5f4HRL7
72Rb0rhInuOchIHxWN1LBixy73gCxluq41mREClFxYtnFlTzbna3XKgfltFqRGKjUjUu4j0dkAKc
SbNGjGIWmq8ZwK47Lzd360JhUv893RmRA1kHTUcHvLrx64QGo1n9O8PN9Mul5ZoolIsbSZtjLfSc
/9fFegobVI7jmSj/jUHffJXEfjTVp//9JKq03aolE7wQWdGVneo4fo5ZZd/2Jnc+VJxBAVVfQUtv
c6been2r2BaDSMHjPBGwfUvXhf5Pg+kK6tZZBmfRXZxqmjD6bF1kSz/ROxT/4c9zVqBpV7TJnko+
vzNRI5E37j6BAn/V59MudoefSwvDMtDXC4DFo6PeVgg/Ts8bPZa51PMsJVkTLVBDlpKH3j7hke3n
Cu9rFz7hWI3Wcv0LsPjyZDJzZuGnRIOC7KWyeztysUSba+zhwy1kVxlMiZRYgzMsyEpOUpdW8ked
YmjTPlDSZKXrfQ8VyeCOV/MoUGm7wj+P0EWzA0Tqffj8eDeChFTBxJwHpRxeLQzb/yUKoJtgrRSK
0QW2b5A4OCGFkwTfjPdAagl8lzm+994EtYkWo9zPj7Jvx2bxYYW/eeUW7xl0kItSpiYBL7uBUIvr
yTkrogY6qO44iHjP8+6o5rxZqhM6iK43caeWV61WJhNVHojv5T/BdmAER4V8eISXEvF2A8QHoRt5
XgN60MZegrcE++oD1zyVgM9+HocV6FBb+PGXJSY4t8gufy3ERndZItf0KB7v21RjGKNmGhPc+cUW
REEItwTZv+g6humbqOHO7kI6utjVnF3RfjookKnI0RVWCWSI/73HMgPEZdmt19wul9UMJJtIFYgI
3l61O2YNaye9OPC6kowPsQ+yC6zUZspvY8PvQqUQnjZ2/3kqU71wJ8MlcDr5FA4EUTYCjhmibW52
lhMMZoFUfBtUMRjb5xiDHvezl1KQ354/QdvO3YewX7USRw9DTGvmIZ6uDazhFgxYGGbXQuPTQ4fB
SRgMcm/dbTnBZYrQkCuOhP58BwdkbzU2PAh1d95ZnTrfp/pZLkUXpjOGIRdtDxT7vcOpDnsK8zW3
2GIMjjiE2h8S5k5eVpXG7hLPqS8AdeBWHg4az4AO/uSj8m+jtU6gVQ07lO2XB8zJrHCsvUM+y0tj
ebQNmJHTWxMbl3xSdMyCiniyjrNTSUCYpp9BQxlyvshX8iCeaofRQt0FOThLx1NFNbkaI5Z9/q1/
scttEflrRUPgqkGT95wxdXzN2w6s6TUya/3a2Ncw6M9IGWffw3L9E7yRRhNvwLgbbgf8l2i1scA+
BZSDpMHDMF8x4p4VWYKDSmk4IKaaH9zQ7oYkvAysli6+v0dgOro8JDKLTcYalrYR57OjdHXMvDKW
HTTMpSAWczcVJa30G8/g7Nwd0/kzIutnw8i/UyJcQMgaUbyQLbg9jXefdIuCFkHIOXslYEtMKtlh
oB93WzRwk8kiHNaKyuO6MqckBGD0C2ac8+exjisWotbdrZsrAgbtyIHllbXQWj1s6Hkhw9AuTEUu
0ee7EWw/BAQsS340Im8vWi5WqaTiMmsf0PkQ9B3/GKGGSium0fWEjZloO9GFFj0SMPS3uKd53d8n
iHhm8gT5oHwE5ERZfgV2Y/PvWetXhQxq+Q8u4gMtCoIsY1bEZuf0sgEOLgIXNBA+u1doSuOVs5bk
ffrbckEkuUlc2DVkEP9JQLcVNGOzw3sHjbw8IrVedBZMrxKCqhsWuYfrjQjrpTe9+BZwTlpJspJB
9XLJH/vysmmFUzZvqFRJR9OK3BtnJi/45u4dz0ovQCBtb5LpxJ8a1xsKBrRt7v8xYrUra0VirpM0
vnSR43eKVaVkGceSNIOcRm31C41+YeAdQoB6aOm1fQOKjGaJ5HLpodGbIi78dsItPbgkW4N8fzde
B7K9TXitHRZ6Fs8dOgAQO0H9QnDaHboWGpkW4EZ/2hX6+Y87+haU5bEyNwHTIR5MEKghEDc0Lu/8
MabkiZM4hTOBcq7yCw471byaU5HIcKnoaQI6SnGR2SQiFTbkQBgLPOhke3qioXcD5OQ2UG1hDwBc
3pcUowFg1iijF30q5ckyxV3X2yrBgGOQv2xaKS+e9irK0CCC/eptdKntzWuenFWyI17QKJx/Cd7c
OzrDLHacl2VY8k/96wVgNSeJQzR33QikqpX7u6XnVfFEaatkez7EoRUoorEh3GJ8aBZ6avHQNKUP
rITo3FNKeURkKaefhjk2tT0xJ5vhCzP5TYLC44oINAIjOwzPuY+es+sTcS6IOIWlIEqYt7tJeCHL
IuNMGiellY+z/RqS1uPLQp7u7/OOWygwsECfNdcHcisgGpP7jJ9DYv4eku0ji/sZwnIK53IKcg1N
fdj45hZGAKmhXu8crVMdl89cko6VBaMX82b4B1f5sCImjKVuWjs7ggjAvlMH7ZZB+186F7HLA25D
47pFZC/q5DO+2zkXd89EcMj0wGkJjIzAdUZesXZLsoB+sChZcQTFwieXzpaXBKRGwdxKhoFOMuqn
NY7Eq38ujFosaruS6QQLJYaV1ZKPpI30omzpW0uHpm//eGCOOm1A5NQzHg9BdQqyffEbzjrIf9e/
AhJU6QUCSKR10d44V3mMsqssJ6KzSN0N4ghEGYF0WuvKDsbmPXsgvPW/njTozWN0D6mQUlLVdMRW
BQf9l7O8A0dhLLbMMalCLT3dgD87AHbbrp+b4dWZoP3uVvnEsA5RWvdYGhDy
`pragma protect end_protected
