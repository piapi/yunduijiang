
`timescale 1 ns / 1 ps

module rgmii_rx(
//    input              idelay_clk  , //200Mhz时钟，IDELAY时钟
    
    //以太网RGMII接口
    input              rgmii_rxc   , //RGMII接收时钟
    input              rgmii_rx_ctl, //RGMII接收数据控制信号
    input       [3:0]  rgmii_rxd   , //RGMII接收数据    

    //以太网GMII接口
    output             gmii_rx_clk , //GMII接收时钟
    output             gmii_rx_dv  , //GMII接收数据有效信号
    output      [7:0]  gmii_rxd      //GMII接收数据   
    );

//parameter define
//parameter IDELAY_VALUE = 0;
parameter  DELAY_VALUE=50;//;0~127

//wire define
wire         rgmii_rxc_bufg;     //全局时钟缓存
wire         rgmii_rxc_bufio;    //全局时钟IO缓存
wire  [3:0]  rgmii_rxd_delay;    //rgmii_rxd输入延时
wire         rgmii_rx_ctl_delay; //rgmii_rx_ctl输入延时
wire  [1:0]  gmii_rxdv_t;        //两位GMII接收有效信号 

//*****************************************************
//**                    main code
//*****************************************************

assign gmii_rx_clk = rgmii_rxc_bufg;
assign gmii_rx_dv = gmii_rxdv_t[0] & gmii_rxdv_t[1];

//全局时钟缓存
BUFG BUFG_inst (
  .I            (rgmii_rxc),     // 1-bit input: Clock input
  .O            (rgmii_rxc_bufg) // 1-bit output: Clock output
);

//全局时钟IO缓存
BUFG BUFIO_inst_1 (
  .I            (rgmii_rxc),      // 1-bit input: Clock input
  .O            (rgmii_rxc_bufio) // 1-bit output: Clock output
);

//输入延时控制
// Specifies group name for associated IDELAYs/ODELAYs and IDELAYCTRL
//(* IODELAY_GROUP = "rgmii_rx_delay" *) 
//IDELAYCTRL  IDELAYCTRL_inst (
//    .RDY(),                      // 1-bit output: Ready output
//    .REFCLK(idelay_clk),         // 1-bit input: Reference clock input
//    .RST(1'b0)                   // 1-bit input: Active high reset input
//);

//rgmii_rx_ctl输入延时与双沿采样
//(* IODELAY_GROUP = "rgmii_rx_delay" *) 
//IDELAYE2 #(
//  .IDELAY_TYPE     ("FIXED"),           // FIXED, VARIABLE, VAR_LOAD, VAR_LOAD_PIPE
//  .IDELAY_VALUE    (IDELAY_VALUE),      // Input delay tap setting (0-31)
//  .REFCLK_FREQUENCY(200.0)              // IDELAYCTRL clock input frequency in MHz 
//)
//u_delay_rx_ctrl (
//  .CNTVALUEOUT     (),                  // 5-bit output: Counter value output
//  .DATAOUT         (rgmii_rx_ctl_delay),// 1-bit output: Delayed data output
//  .C               (1'b0),              // 1-bit input: Clock input
//  .CE              (1'b0),              // 1-bit input: enable increment/decrement
//  .CINVCTRL        (1'b0),              // 1-bit input: Dynamic clock inversion input
//  .CNTVALUEIN      (5'b0),              // 5-bit input: Counter value input
//  .DATAIN          (1'b0),              // 1-bit input: Internal delay data input
//  .IDATAIN         (rgmii_rx_ctl),      // 1-bit input: Data input from the I/O
//  .INC             (1'b0),              // 1-bit input: Increment / Decrement tap delay
//  .LD              (1'b0),              // 1-bit input: Load IDELAY_VALUE input
//  .LDPIPEEN        (1'b0),              // 1-bit input: Enable PIPELINE register
//  .REGRST          (1'b0)               // 1-bit input: Active-high reset tap-delay input
//);

//输入双沿采样寄存器
//IDDR #(
//    .DDR_CLK_EDGE("SAME_EDGE_PIPELINED"),// "OPPOSITE_EDGE", "SAME_EDGE" 
//                                            or "SAME_EDGE_PIPELINED" 
//    .INIT_Q1  (1'b0),                   // Initial value of Q1: 1'b0 or 1'b1
//    .INIT_Q2  (1'b0),                   // Initial value of Q2: 1'b0 or 1'b1
//    .SRTYPE   ("SYNC")                  // Set/Reset type: "SYNC" or "ASYNC" 
//) u_iddr_rx_ctl (
//    .Q1       (gmii_rxdv_t[0]),         // 1-bit output for positive edge of clock
//    .Q2       (gmii_rxdv_t[1]),         // 1-bit output for negative edge of clock
//    .C        (rgmii_rxc_bufio),        // 1-bit clock input
//    .CE       (1'b1),                   // 1-bit clock enable input
//    .D        (rgmii_rx_ctl_delay),     // 1-bit DDR data input
//    .R        (1'b0),                   // 1-bit reset
//    .S        (1'b0)                    // 1-bit set
//);


IODELAY #(.C_STATIC_DLY(DELAY_VALUE))//integer,0~127
        IODELAY_inst_dv1(
        .DO(rgmii_rx_ctl_delay), 
        .DF(), 
        .DI(rgmii_rx_ctl), 
        .SDTAP(0), 
        .SETN(0), 
        .VALUE(0)
        );

		IDDR	  U_IDDR_dv1
						(.Q0(gmii_rxdv_t[0]), 
						.Q1(gmii_rxdv_t[1]), 
						.D(rgmii_rx_ctl_delay), 
						.CLK(rgmii_rxc_bufio) 
						);


//rgmii_rxd输入延时与双沿采样
//genvar i;
//generate for (i=0; i<4; i=i+1)
//    (* IODELAY_GROUP = "rgmii_rx_delay" *) 
//    begin : rxdata_bus
//        输入延时           
//        (* IODELAY_GROUP = "rgmii_rx_delay" *) 
//        IDELAYE2 #(
//          .IDELAY_TYPE     ("FIXED"),           // FIXED,VARIABLE,VAR_LOAD,VAR_LOAD_PIPE
//          .IDELAY_VALUE    (IDELAY_VALUE),      // Input delay tap setting (0-31)    
//          .REFCLK_FREQUENCY(200.0)              // IDELAYCTRL clock input frequency in MHz
//        )
//        u_delay_rxd (
//          .CNTVALUEOUT     (),                  // 5-bit output: Counter value output
//          .DATAOUT         (rgmii_rxd_delay[i]),// 1-bit output: Delayed data output
//          .C               (1'b0),              // 1-bit input: Clock input
//          .CE              (1'b0),              // 1-bit input: enable increment/decrement
//          .CINVCTRL        (1'b0),              // 1-bit input: Dynamic clock inversion
//          .CNTVALUEIN      (5'b0),              // 5-bit input: Counter value input
//          .DATAIN          (1'b0),              // 1-bit input: Internal delay data input
//          .IDATAIN         (rgmii_rxd[i]),      // 1-bit input: Data input from the I/O
//          .INC             (1'b0),              // 1-bit input: Inc/Decrement tap delay
//          .LD              (1'b0),              // 1-bit input: Load IDELAY_VALUE input
//          .LDPIPEEN        (1'b0),              // 1-bit input: Enable PIPELINE register 
//          .REGRST          (1'b0)               // 1-bit input: Active-high reset tap-delay
//        );
//        
//        输入双沿采样寄存器
//        IDDR #(
//            .DDR_CLK_EDGE("SAME_EDGE_PIPELINED"),// "OPPOSITE_EDGE", "SAME_EDGE" 
//                                                    or "SAME_EDGE_PIPELINED" 
//            .INIT_Q1  (1'b0),                   // Initial value of Q1: 1'b0 or 1'b1
//            .INIT_Q2  (1'b0),                   // Initial value of Q2: 1'b0 or 1'b1
//            .SRTYPE   ("SYNC")                  // Set/Reset type: "SYNC" or "ASYNC" 
//        ) u_iddr_rxd (
//            .Q1       (gmii_rxd[i]),            // 1-bit output for positive edge of clock
//            .Q2       (gmii_rxd[4+i]),          // 1-bit output for negative edge of clock
//            .C        (rgmii_rxc_bufio),        // 1-bit clock input rgmii_rxc_bufio
//            .CE       (1'b1),                   // 1-bit clock enable input
//            .D        (rgmii_rxd_delay[i]),     // 1-bit DDR data input
//            .R        (1'b0),                   // 1-bit reset
//            .S        (1'b0)                    // 1-bit set
//        );
//    end
//endgenerate
   generate
	genvar m ;
		for(m=0;m<=3;m=m+1) 
		begin
                IODELAY #(.C_STATIC_DLY(DELAY_VALUE))//integer,0~127
                IODELAY_inst_dq1(
                .DO(rgmii_rxd_delay[m]), 
                .DF(), 
                .DI(rgmii_rxd[m]), 
                .SDTAP(0), 
                .SETN(0), 
                .VALUE(0)
                );

		end
   endgenerate

   generate
	genvar i ;
		for(i=0;i<=3;i=i+1) 
		begin
		IDDR	  U_IDDR_dq1
						(.Q0(gmii_rxd[i]), 
						.Q1(gmii_rxd[i+4]), 
						.D(rgmii_rxd_delay[i]), 
						.CLK(rgmii_rxc_bufio) 
						);
		end
   endgenerate

endmodule